-- VHDL produced by vc2vhdl from virtual circuit (vc) description 
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;xxxxxxx
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;
library work;
use work.ahir_system_global_package.all;
entity vector_control_daemon is -- 
  generic (tag_length : integer); 
  port ( -- 
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic;
    in_data_pipe_read_req : out  std_logic_vector(0 downto 0);
    in_data_pipe_read_ack : in   std_logic_vector(0 downto 0);
    in_data_pipe_read_data : in   std_logic_vector(31 downto 0);
    out_data_pipe_write_req : out  std_logic_vector(0 downto 0);
    out_data_pipe_write_ack : in   std_logic_vector(0 downto 0);
    out_data_pipe_write_data : out  std_logic_vector(31 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) -- 
  );
  -- 
end entity vector_control_daemon;
architecture Default of vector_control_daemon is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal default_zero_sig: std_logic;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal vector_control_daemon_CP_10259_start: Boolean;
  signal vector_control_daemon_CP_10259_symbol: Boolean;
  -- links between control-path and data-path
  signal RPIPE_in_data_2071_inst_req_1 : boolean;
  signal RPIPE_in_data_2071_inst_ack_1 : boolean;
  signal ADD_f32_f32_2093_inst_req_0 : boolean;
  signal ADD_f32_f32_2093_inst_ack_0 : boolean;
  signal RPIPE_in_data_2068_inst_req_0 : boolean;
  signal RPIPE_in_data_2068_inst_ack_0 : boolean;
  signal RPIPE_in_data_2077_inst_ack_1 : boolean;
  signal UGT_u32_u1_2394_inst_req_0 : boolean;
  signal MUL_f32_f32_2099_inst_req_0 : boolean;
  signal MUL_f32_f32_2099_inst_ack_0 : boolean;
  signal MUL_f32_f32_2099_inst_req_1 : boolean;
  signal MUL_f32_f32_2099_inst_ack_1 : boolean;
  signal RPIPE_in_data_2077_inst_req_0 : boolean;
  signal RPIPE_in_data_2077_inst_ack_0 : boolean;
  signal RPIPE_in_data_2077_inst_req_1 : boolean;
  signal if_stmt_2437_branch_ack_1 : boolean;
  signal type_cast_2104_inst_req_0 : boolean;
  signal type_cast_2104_inst_ack_0 : boolean;
  signal type_cast_2104_inst_req_1 : boolean;
  signal UGT_u32_u1_2394_inst_ack_0 : boolean;
  signal RPIPE_in_data_2074_inst_req_1 : boolean;
  signal RPIPE_in_data_2074_inst_ack_1 : boolean;
  signal MUL_f32_f32_2088_inst_req_1 : boolean;
  signal MUL_f32_f32_2088_inst_ack_1 : boolean;
  signal SHL_u32_u32_2354_inst_ack_1 : boolean;
  signal MUL_f32_f32_2088_inst_req_0 : boolean;
  signal MUL_f32_f32_2088_inst_ack_0 : boolean;
  signal RPIPE_in_data_2068_inst_req_1 : boolean;
  signal RPIPE_in_data_2068_inst_ack_1 : boolean;
  signal AND_u32_u32_3460_inst_ack_1 : boolean;
  signal AND_u32_u32_3460_inst_req_1 : boolean;
  signal SLT_f64_u1_2110_inst_ack_1 : boolean;
  signal RPIPE_in_data_2071_inst_req_0 : boolean;
  signal RPIPE_in_data_2071_inst_ack_0 : boolean;
  signal if_stmt_2437_branch_req_0 : boolean;
  signal type_cast_2104_inst_ack_1 : boolean;
  signal SLT_f64_u1_2110_inst_req_0 : boolean;
  signal SLT_f64_u1_2110_inst_ack_0 : boolean;
  signal SLT_f64_u1_2110_inst_req_1 : boolean;
  signal RPIPE_in_data_2074_inst_req_0 : boolean;
  signal RPIPE_in_data_2074_inst_ack_0 : boolean;
  signal LSHR_u32_u32_2388_inst_ack_1 : boolean;
  signal SHL_u32_u32_2354_inst_ack_0 : boolean;
  signal LSHR_u32_u32_2388_inst_req_1 : boolean;
  signal SUB_f32_f32_2082_inst_req_0 : boolean;
  signal SUB_f32_f32_2082_inst_ack_0 : boolean;
  signal SUB_f32_f32_2082_inst_req_1 : boolean;
  signal SUB_f32_f32_2082_inst_ack_1 : boolean;
  signal ADD_f32_f32_2093_inst_req_1 : boolean;
  signal ADD_f32_f32_2093_inst_ack_1 : boolean;
  signal UGT_u32_u1_2394_inst_req_1 : boolean;
  signal UGT_u32_u1_2394_inst_ack_1 : boolean;
  signal if_stmt_2396_branch_req_0 : boolean;
  signal if_stmt_2396_branch_ack_1 : boolean;
  signal if_stmt_2396_branch_ack_0 : boolean;
  signal SHL_u32_u32_2424_inst_req_0 : boolean;
  signal if_stmt_2112_branch_req_0 : boolean;
  signal if_stmt_2112_branch_ack_1 : boolean;
  signal if_stmt_2112_branch_ack_0 : boolean;
  signal SGT_f64_u1_2123_inst_req_0 : boolean;
  signal SGT_f64_u1_2123_inst_ack_0 : boolean;
  signal SGT_f64_u1_2123_inst_req_1 : boolean;
  signal SGT_f64_u1_2123_inst_ack_1 : boolean;
  signal if_stmt_2125_branch_req_0 : boolean;
  signal if_stmt_2125_branch_ack_1 : boolean;
  signal if_stmt_2125_branch_ack_0 : boolean;
  signal MUL_f32_f32_2149_inst_req_0 : boolean;
  signal MUL_f32_f32_2149_inst_ack_0 : boolean;
  signal MUL_f32_f32_2149_inst_req_1 : boolean;
  signal MUL_f32_f32_2149_inst_ack_1 : boolean;
  signal ADD_f32_f32_2154_inst_req_0 : boolean;
  signal ADD_f32_f32_2154_inst_ack_0 : boolean;
  signal ADD_f32_f32_2154_inst_req_1 : boolean;
  signal ADD_f32_f32_2154_inst_ack_1 : boolean;
  signal SLT_f32_u1_2160_inst_req_0 : boolean;
  signal SLT_f32_u1_2160_inst_ack_0 : boolean;
  signal SLT_f32_u1_2160_inst_req_1 : boolean;
  signal SLT_f32_u1_2160_inst_ack_1 : boolean;
  signal if_stmt_2162_branch_req_0 : boolean;
  signal if_stmt_2162_branch_ack_1 : boolean;
  signal if_stmt_2162_branch_ack_0 : boolean;
  signal SGT_f32_u1_2173_inst_req_0 : boolean;
  signal SGT_f32_u1_2173_inst_ack_0 : boolean;
  signal SGT_f32_u1_2173_inst_req_1 : boolean;
  signal SGT_f32_u1_2173_inst_ack_1 : boolean;
  signal if_stmt_2437_branch_ack_0 : boolean;
  signal SHL_u32_u32_2354_inst_req_0 : boolean;
  signal if_stmt_2175_branch_req_0 : boolean;
  signal if_stmt_2175_branch_ack_1 : boolean;
  signal if_stmt_2175_branch_ack_0 : boolean;
  signal LSHR_u32_u32_2388_inst_ack_0 : boolean;
  signal LSHR_u32_u32_2388_inst_req_0 : boolean;
  signal MUL_f32_f32_2186_inst_req_0 : boolean;
  signal MUL_f32_f32_2186_inst_ack_0 : boolean;
  signal MUL_f32_f32_2186_inst_req_1 : boolean;
  signal MUL_f32_f32_2186_inst_ack_1 : boolean;
  signal SHL_u32_u32_2430_inst_ack_0 : boolean;
  signal ULT_u32_u1_2435_inst_ack_0 : boolean;
  signal ULT_u32_u1_2435_inst_ack_1 : boolean;
  signal ULT_u32_u1_2435_inst_req_1 : boolean;
  signal type_cast_2203_inst_req_0 : boolean;
  signal type_cast_2203_inst_ack_0 : boolean;
  signal type_cast_2203_inst_req_1 : boolean;
  signal type_cast_2203_inst_ack_1 : boolean;
  signal SHL_u32_u32_2430_inst_req_0 : boolean;
  signal SHL_u32_u32_2430_inst_ack_1 : boolean;
  signal SGT_f64_u1_2209_inst_req_0 : boolean;
  signal SGT_f64_u1_2209_inst_ack_0 : boolean;
  signal OR_u32_u32_2366_inst_ack_1 : boolean;
  signal SGT_f64_u1_2209_inst_req_1 : boolean;
  signal SGT_f64_u1_2209_inst_ack_1 : boolean;
  signal SHL_u32_u32_2424_inst_ack_0 : boolean;
  signal OR_u32_u32_2366_inst_req_1 : boolean;
  signal LSHR_u32_u32_2728_inst_req_0 : boolean;
  signal MUL_f32_f32_2695_inst_ack_0 : boolean;
  signal if_stmt_2211_branch_req_0 : boolean;
  signal ULT_u32_u1_2435_inst_req_0 : boolean;
  signal if_stmt_2211_branch_ack_1 : boolean;
  signal if_stmt_2211_branch_ack_0 : boolean;
  signal OR_u32_u32_2366_inst_ack_0 : boolean;
  signal OR_u32_u32_2366_inst_req_0 : boolean;
  signal SHL_u32_u32_2430_inst_req_1 : boolean;
  signal SGT_f64_u1_2222_inst_req_0 : boolean;
  signal SGT_f64_u1_2222_inst_ack_0 : boolean;
  signal SGT_f64_u1_2222_inst_req_1 : boolean;
  signal SGT_f64_u1_2222_inst_ack_1 : boolean;
  signal SHL_u32_u32_2354_inst_req_1 : boolean;
  signal if_stmt_2343_branch_ack_0 : boolean;
  signal if_stmt_2224_branch_req_0 : boolean;
  signal if_stmt_2224_branch_ack_1 : boolean;
  signal if_stmt_2224_branch_ack_0 : boolean;
  signal if_stmt_2343_branch_ack_1 : boolean;
  signal MUL_f32_f32_2235_inst_req_0 : boolean;
  signal MUL_f32_f32_2235_inst_ack_0 : boolean;
  signal MUL_f32_f32_2235_inst_req_1 : boolean;
  signal MUL_f32_f32_2235_inst_ack_1 : boolean;
  signal AND_u32_u32_2360_inst_ack_1 : boolean;
  signal AND_u32_u32_2360_inst_req_1 : boolean;
  signal ADD_f32_f32_2241_inst_req_0 : boolean;
  signal ADD_f32_f32_2241_inst_ack_0 : boolean;
  signal ADD_f32_f32_2241_inst_req_1 : boolean;
  signal ADD_f32_f32_2241_inst_ack_1 : boolean;
  signal AND_u32_u32_2360_inst_ack_0 : boolean;
  signal AND_u32_u32_2360_inst_req_0 : boolean;
  signal MUL_f32_f32_2247_inst_req_0 : boolean;
  signal MUL_f32_f32_2247_inst_ack_0 : boolean;
  signal MUL_f32_f32_2247_inst_req_1 : boolean;
  signal MUL_f32_f32_2247_inst_ack_1 : boolean;
  signal SHL_u32_u32_2424_inst_ack_1 : boolean;
  signal SHL_u32_u32_2424_inst_req_1 : boolean;
  signal SGT_f64_u1_2255_inst_req_0 : boolean;
  signal SGT_f64_u1_2255_inst_ack_0 : boolean;
  signal SGT_f64_u1_2255_inst_req_1 : boolean;
  signal SGT_f64_u1_2255_inst_ack_1 : boolean;
  signal if_stmt_2257_branch_req_0 : boolean;
  signal LSHR_u32_u32_2728_inst_ack_0 : boolean;
  signal LSHR_u32_u32_2740_inst_req_0 : boolean;
  signal if_stmt_2257_branch_ack_1 : boolean;
  signal if_stmt_2257_branch_ack_0 : boolean;
  signal MUL_f32_f32_2268_inst_req_0 : boolean;
  signal MUL_f32_f32_2268_inst_ack_0 : boolean;
  signal MUL_f32_f32_2268_inst_req_1 : boolean;
  signal MUL_f32_f32_2268_inst_ack_1 : boolean;
  signal ADD_f32_f32_2274_inst_req_0 : boolean;
  signal ADD_f32_f32_2274_inst_ack_0 : boolean;
  signal ADD_f32_f32_2274_inst_req_1 : boolean;
  signal ADD_f32_f32_2274_inst_ack_1 : boolean;
  signal NEQ_i32_u1_3028_inst_ack_0 : boolean;
  signal MUL_f32_f32_2280_inst_req_0 : boolean;
  signal MUL_f32_f32_2280_inst_ack_0 : boolean;
  signal MUL_f32_f32_2280_inst_req_1 : boolean;
  signal MUL_f32_f32_2280_inst_ack_1 : boolean;
  signal EQ_f32_u1_2715_inst_req_0 : boolean;
  signal EQ_f32_u1_2715_inst_ack_0 : boolean;
  signal MUL_f32_f32_2288_inst_req_0 : boolean;
  signal MUL_f32_f32_2288_inst_ack_0 : boolean;
  signal MUL_f32_f32_2695_inst_ack_1 : boolean;
  signal MUL_f32_f32_2288_inst_req_1 : boolean;
  signal MUL_f32_f32_2288_inst_ack_1 : boolean;
  signal LSHR_u32_u32_2740_inst_ack_1 : boolean;
  signal EQ_f32_u1_2715_inst_req_1 : boolean;
  signal ADD_f32_f32_2294_inst_req_0 : boolean;
  signal ADD_f32_f32_2294_inst_ack_0 : boolean;
  signal ADD_f32_f32_2294_inst_req_1 : boolean;
  signal ADD_f32_f32_2294_inst_ack_1 : boolean;
  signal EQ_f32_u1_2715_inst_ack_1 : boolean;
  signal MUL_f32_f32_2300_inst_req_0 : boolean;
  signal MUL_f32_f32_2300_inst_ack_0 : boolean;
  signal MUL_f32_f32_2695_inst_req_0 : boolean;
  signal MUL_f32_f32_2300_inst_req_1 : boolean;
  signal MUL_f32_f32_2300_inst_ack_1 : boolean;
  signal MUL_f32_f32_2320_inst_req_0 : boolean;
  signal MUL_f32_f32_2320_inst_ack_0 : boolean;
  signal MUL_f32_f32_2320_inst_req_1 : boolean;
  signal MUL_f32_f32_2320_inst_ack_1 : boolean;
  signal MUL_f32_f32_2326_inst_req_0 : boolean;
  signal MUL_f32_f32_2326_inst_ack_0 : boolean;
  signal MUL_f32_f32_2326_inst_req_1 : boolean;
  signal MUL_f32_f32_2326_inst_ack_1 : boolean;
  signal ADD_f32_f32_2331_inst_req_0 : boolean;
  signal ADD_f32_f32_2331_inst_ack_0 : boolean;
  signal ADD_f32_f32_2331_inst_req_1 : boolean;
  signal ADD_f32_f32_2331_inst_ack_1 : boolean;
  signal type_cast_2335_inst_req_0 : boolean;
  signal type_cast_2335_inst_ack_0 : boolean;
  signal type_cast_2335_inst_req_1 : boolean;
  signal type_cast_2335_inst_ack_1 : boolean;
  signal EQ_f32_u1_2341_inst_req_0 : boolean;
  signal EQ_f32_u1_2341_inst_ack_0 : boolean;
  signal EQ_f32_u1_2341_inst_req_1 : boolean;
  signal EQ_f32_u1_2341_inst_ack_1 : boolean;
  signal if_stmt_2343_branch_req_0 : boolean;
  signal ADD_u32_u32_2473_inst_req_0 : boolean;
  signal ADD_u32_u32_2473_inst_ack_0 : boolean;
  signal ADD_u32_u32_2473_inst_req_1 : boolean;
  signal ADD_u32_u32_2473_inst_ack_1 : boolean;
  signal SUB_u32_u32_2478_inst_req_0 : boolean;
  signal SUB_u32_u32_2478_inst_ack_0 : boolean;
  signal SUB_u32_u32_2478_inst_req_1 : boolean;
  signal SUB_u32_u32_2478_inst_ack_1 : boolean;
  signal ULT_u32_u1_2484_inst_req_0 : boolean;
  signal ULT_u32_u1_2484_inst_ack_0 : boolean;
  signal ULT_u32_u1_2484_inst_req_1 : boolean;
  signal ULT_u32_u1_2484_inst_ack_1 : boolean;
  signal if_stmt_2486_branch_req_0 : boolean;
  signal if_stmt_2486_branch_ack_1 : boolean;
  signal if_stmt_2486_branch_ack_0 : boolean;
  signal LSHR_u32_u32_2502_inst_req_0 : boolean;
  signal LSHR_u32_u32_2502_inst_ack_0 : boolean;
  signal LSHR_u32_u32_2502_inst_req_1 : boolean;
  signal LSHR_u32_u32_2502_inst_ack_1 : boolean;
  signal AND_u32_u32_2508_inst_req_0 : boolean;
  signal AND_u32_u32_2508_inst_ack_0 : boolean;
  signal AND_u32_u32_2508_inst_req_1 : boolean;
  signal AND_u32_u32_2508_inst_ack_1 : boolean;
  signal AND_u32_u32_2514_inst_req_0 : boolean;
  signal AND_u32_u32_2514_inst_ack_0 : boolean;
  signal AND_u32_u32_2514_inst_req_1 : boolean;
  signal AND_u32_u32_2514_inst_ack_1 : boolean;
  signal ADD_u32_u32_2520_inst_req_0 : boolean;
  signal ADD_u32_u32_2520_inst_ack_0 : boolean;
  signal ADD_u32_u32_2520_inst_req_1 : boolean;
  signal ADD_u32_u32_2520_inst_ack_1 : boolean;
  signal AND_u32_u32_2526_inst_req_0 : boolean;
  signal AND_u32_u32_2526_inst_ack_0 : boolean;
  signal AND_u32_u32_2526_inst_req_1 : boolean;
  signal AND_u32_u32_2526_inst_ack_1 : boolean;
  signal EQ_u32_u1_2532_inst_req_0 : boolean;
  signal EQ_u32_u1_2532_inst_ack_0 : boolean;
  signal EQ_u32_u1_2532_inst_req_1 : boolean;
  signal EQ_u32_u1_2532_inst_ack_1 : boolean;
  signal type_cast_2536_inst_req_0 : boolean;
  signal type_cast_2536_inst_ack_0 : boolean;
  signal type_cast_2536_inst_req_1 : boolean;
  signal type_cast_2536_inst_ack_1 : boolean;
  signal AND_u32_u32_2734_inst_ack_1 : boolean;
  signal OR_u32_u32_2764_inst_ack_1 : boolean;
  signal NEQ_i32_u1_2540_inst_req_0 : boolean;
  signal NEQ_i32_u1_2540_inst_ack_0 : boolean;
  signal NEQ_i32_u1_2540_inst_req_1 : boolean;
  signal NEQ_i32_u1_2540_inst_ack_1 : boolean;
  signal AND_u32_u32_2734_inst_req_1 : boolean;
  signal OR_u32_u32_2764_inst_req_1 : boolean;
  signal SHL_u32_u32_2752_inst_ack_1 : boolean;
  signal type_cast_2709_inst_ack_1 : boolean;
  signal LSHR_u32_u32_2740_inst_req_1 : boolean;
  signal SHL_u32_u32_2752_inst_req_1 : boolean;
  signal type_cast_2709_inst_req_1 : boolean;
  signal SHL_u32_u32_2752_inst_ack_0 : boolean;
  signal SHL_u32_u32_2752_inst_req_0 : boolean;
  signal AND_u1_u1_2545_inst_req_0 : boolean;
  signal AND_u1_u1_2545_inst_ack_0 : boolean;
  signal AND_u1_u1_2545_inst_req_1 : boolean;
  signal AND_u1_u1_2545_inst_ack_1 : boolean;
  signal OR_u32_u32_2764_inst_ack_0 : boolean;
  signal NEQ_i32_u1_3028_inst_req_1 : boolean;
  signal if_stmt_2717_branch_req_0 : boolean;
  signal type_cast_2709_inst_ack_0 : boolean;
  signal type_cast_2679_inst_ack_1 : boolean;
  signal type_cast_2709_inst_req_0 : boolean;
  signal if_stmt_2547_branch_req_0 : boolean;
  signal type_cast_2679_inst_req_1 : boolean;
  signal if_stmt_2547_branch_ack_1 : boolean;
  signal if_stmt_2547_branch_ack_0 : boolean;
  signal SHL_u32_u32_2574_inst_req_0 : boolean;
  signal SHL_u32_u32_2574_inst_ack_0 : boolean;
  signal MUL_f32_f32_2695_inst_req_1 : boolean;
  signal SHL_u32_u32_2574_inst_req_1 : boolean;
  signal SHL_u32_u32_2574_inst_ack_1 : boolean;
  signal OR_u32_u32_2764_inst_req_0 : boolean;
  signal AND_u32_u32_2580_inst_req_0 : boolean;
  signal AND_u32_u32_2580_inst_ack_0 : boolean;
  signal AND_u32_u32_2580_inst_req_1 : boolean;
  signal AND_u32_u32_2580_inst_ack_1 : boolean;
  signal type_cast_2705_inst_ack_1 : boolean;
  signal type_cast_2705_inst_req_1 : boolean;
  signal EQ_u32_u1_2586_inst_req_0 : boolean;
  signal EQ_u32_u1_2586_inst_ack_0 : boolean;
  signal EQ_u32_u1_2586_inst_req_1 : boolean;
  signal EQ_u32_u1_2586_inst_ack_1 : boolean;
  signal AND_u32_u32_2734_inst_ack_0 : boolean;
  signal AND_u32_u32_2746_inst_ack_1 : boolean;
  signal AND_u32_u32_2746_inst_req_1 : boolean;
  signal type_cast_2705_inst_ack_0 : boolean;
  signal type_cast_2705_inst_req_0 : boolean;
  signal LSHR_u32_u32_2740_inst_ack_0 : boolean;
  signal type_cast_2590_inst_req_0 : boolean;
  signal type_cast_2590_inst_ack_0 : boolean;
  signal type_cast_2590_inst_req_1 : boolean;
  signal type_cast_2590_inst_ack_1 : boolean;
  signal AND_u32_u32_2734_inst_req_0 : boolean;
  signal AND_u32_u32_2746_inst_ack_0 : boolean;
  signal AND_u32_u32_2746_inst_req_0 : boolean;
  signal NEQ_i32_u1_2594_inst_req_0 : boolean;
  signal NEQ_i32_u1_2594_inst_ack_0 : boolean;
  signal NEQ_i32_u1_2594_inst_req_1 : boolean;
  signal NEQ_i32_u1_2594_inst_ack_1 : boolean;
  signal AND_u32_u32_2758_inst_req_1 : boolean;
  signal AND_u32_u32_2758_inst_ack_1 : boolean;
  signal LSHR_u32_u32_2728_inst_ack_1 : boolean;
  signal LSHR_u32_u32_2728_inst_req_1 : boolean;
  signal MUL_f32_f32_2701_inst_ack_1 : boolean;
  signal AND_u1_u1_2599_inst_req_0 : boolean;
  signal AND_u1_u1_2599_inst_ack_0 : boolean;
  signal MUL_f32_f32_2701_inst_req_1 : boolean;
  signal AND_u1_u1_2599_inst_req_1 : boolean;
  signal AND_u1_u1_2599_inst_ack_1 : boolean;
  signal if_stmt_2717_branch_ack_0 : boolean;
  signal MUL_f32_f32_2701_inst_ack_0 : boolean;
  signal ADD_u32_u32_2605_inst_req_0 : boolean;
  signal ADD_u32_u32_2605_inst_ack_0 : boolean;
  signal MUL_f32_f32_2701_inst_req_0 : boolean;
  signal ADD_u32_u32_2605_inst_req_1 : boolean;
  signal ADD_u32_u32_2605_inst_ack_1 : boolean;
  signal if_stmt_2717_branch_ack_1 : boolean;
  signal type_cast_2679_inst_ack_0 : boolean;
  signal type_cast_2679_inst_req_0 : boolean;
  signal if_stmt_2607_branch_req_0 : boolean;
  signal if_stmt_2607_branch_ack_1 : boolean;
  signal if_stmt_2607_branch_ack_0 : boolean;
  signal ADD_u32_u32_2627_inst_req_0 : boolean;
  signal ADD_u32_u32_2627_inst_ack_0 : boolean;
  signal ADD_u32_u32_2627_inst_req_1 : boolean;
  signal ADD_u32_u32_2627_inst_ack_1 : boolean;
  signal AND_u32_u32_2758_inst_req_0 : boolean;
  signal AND_u32_u32_2758_inst_ack_0 : boolean;
  signal SUB_u32_u32_2632_inst_req_0 : boolean;
  signal SUB_u32_u32_2632_inst_ack_0 : boolean;
  signal SUB_u32_u32_2632_inst_req_1 : boolean;
  signal SUB_u32_u32_2632_inst_ack_1 : boolean;
  signal type_cast_3024_inst_req_0 : boolean;
  signal AND_u32_u32_2653_inst_req_0 : boolean;
  signal AND_u32_u32_2653_inst_ack_0 : boolean;
  signal AND_u32_u32_2653_inst_req_1 : boolean;
  signal AND_u32_u32_2653_inst_ack_1 : boolean;
  signal SHL_u32_u32_2659_inst_req_0 : boolean;
  signal SHL_u32_u32_2659_inst_ack_0 : boolean;
  signal SHL_u32_u32_2659_inst_req_1 : boolean;
  signal SHL_u32_u32_2659_inst_ack_1 : boolean;
  signal NEQ_i32_u1_3028_inst_req_0 : boolean;
  signal type_cast_3024_inst_ack_0 : boolean;
  signal ADD_u32_u32_3061_inst_ack_0 : boolean;
  signal ADD_u32_u32_2665_inst_req_0 : boolean;
  signal ADD_u32_u32_2665_inst_ack_0 : boolean;
  signal ADD_u32_u32_2665_inst_req_1 : boolean;
  signal ADD_u32_u32_2665_inst_ack_1 : boolean;
  signal OR_u32_u32_2670_inst_req_0 : boolean;
  signal OR_u32_u32_2670_inst_ack_0 : boolean;
  signal OR_u32_u32_2670_inst_req_1 : boolean;
  signal OR_u32_u32_2670_inst_ack_1 : boolean;
  signal OR_u32_u32_2675_inst_req_0 : boolean;
  signal OR_u32_u32_2675_inst_ack_0 : boolean;
  signal OR_u32_u32_2675_inst_req_1 : boolean;
  signal OR_u32_u32_2675_inst_ack_1 : boolean;
  signal LSHR_u32_u32_2770_inst_req_0 : boolean;
  signal LSHR_u32_u32_2770_inst_ack_0 : boolean;
  signal LSHR_u32_u32_2770_inst_req_1 : boolean;
  signal LSHR_u32_u32_2770_inst_ack_1 : boolean;
  signal AND_u32_u32_2776_inst_req_0 : boolean;
  signal AND_u32_u32_2776_inst_ack_0 : boolean;
  signal AND_u32_u32_2776_inst_req_1 : boolean;
  signal AND_u32_u32_2776_inst_ack_1 : boolean;
  signal OR_u32_u32_2782_inst_req_0 : boolean;
  signal OR_u32_u32_2782_inst_ack_0 : boolean;
  signal OR_u32_u32_2782_inst_req_1 : boolean;
  signal OR_u32_u32_2782_inst_ack_1 : boolean;
  signal XOR_u32_u32_2787_inst_req_0 : boolean;
  signal XOR_u32_u32_2787_inst_ack_0 : boolean;
  signal XOR_u32_u32_2787_inst_req_1 : boolean;
  signal XOR_u32_u32_2787_inst_ack_1 : boolean;
  signal AND_u32_u32_2793_inst_req_0 : boolean;
  signal AND_u32_u32_2793_inst_ack_0 : boolean;
  signal AND_u32_u32_2793_inst_req_1 : boolean;
  signal AND_u32_u32_2793_inst_ack_1 : boolean;
  signal SUB_u32_u32_2798_inst_req_0 : boolean;
  signal SUB_u32_u32_2798_inst_ack_0 : boolean;
  signal SUB_u32_u32_2798_inst_req_1 : boolean;
  signal SUB_u32_u32_2798_inst_ack_1 : boolean;
  signal switch_stmt_2800_branch_default_req_0 : boolean;
  signal switch_stmt_2800_select_expr_0_req_0 : boolean;
  signal switch_stmt_2800_select_expr_0_ack_0 : boolean;
  signal switch_stmt_2800_select_expr_0_req_1 : boolean;
  signal switch_stmt_2800_select_expr_0_ack_1 : boolean;
  signal switch_stmt_2800_branch_0_req_0 : boolean;
  signal switch_stmt_2800_select_expr_1_req_0 : boolean;
  signal switch_stmt_2800_select_expr_1_ack_0 : boolean;
  signal switch_stmt_2800_select_expr_1_req_1 : boolean;
  signal switch_stmt_2800_select_expr_1_ack_1 : boolean;
  signal switch_stmt_2800_branch_1_req_0 : boolean;
  signal switch_stmt_2800_branch_0_ack_1 : boolean;
  signal switch_stmt_2800_branch_1_ack_1 : boolean;
  signal switch_stmt_2800_branch_default_ack_0 : boolean;
  signal LSHR_u32_u32_2831_inst_req_0 : boolean;
  signal LSHR_u32_u32_2831_inst_ack_0 : boolean;
  signal LSHR_u32_u32_2831_inst_req_1 : boolean;
  signal LSHR_u32_u32_2831_inst_ack_1 : boolean;
  signal UGT_u32_u1_2836_inst_req_0 : boolean;
  signal UGT_u32_u1_2836_inst_ack_0 : boolean;
  signal UGT_u32_u1_2836_inst_req_1 : boolean;
  signal UGT_u32_u1_2836_inst_ack_1 : boolean;
  signal if_stmt_2838_branch_req_0 : boolean;
  signal OR_u32_u32_3109_inst_req_1 : boolean;
  signal if_stmt_2838_branch_ack_1 : boolean;
  signal if_stmt_2838_branch_ack_0 : boolean;
  signal SHL_u32_u32_3098_inst_ack_0 : boolean;
  signal SHL_u32_u32_3098_inst_req_0 : boolean;
  signal OR_u32_u32_3109_inst_ack_0 : boolean;
  signal OR_u32_u32_3109_inst_req_0 : boolean;
  signal AND_u32_u32_3092_inst_req_1 : boolean;
  signal SHL_u32_u32_2865_inst_req_0 : boolean;
  signal SHL_u32_u32_2865_inst_ack_0 : boolean;
  signal SHL_u32_u32_2865_inst_req_1 : boolean;
  signal SHL_u32_u32_2865_inst_ack_1 : boolean;
  signal OR_u32_u32_3114_inst_req_1 : boolean;
  signal OR_u32_u32_3114_inst_ack_1 : boolean;
  signal if_stmt_3041_branch_ack_0 : boolean;
  signal SUB_u32_u32_3071_inst_ack_0 : boolean;
  signal type_cast_3024_inst_ack_1 : boolean;
  signal SHL_u32_u32_2871_inst_req_0 : boolean;
  signal SHL_u32_u32_2871_inst_ack_0 : boolean;
  signal SHL_u32_u32_2871_inst_req_1 : boolean;
  signal SHL_u32_u32_2871_inst_ack_1 : boolean;
  signal AND_u32_u32_3460_inst_ack_0 : boolean;
  signal if_stmt_3041_branch_ack_1 : boolean;
  signal AND_u32_u32_3092_inst_ack_0 : boolean;
  signal if_stmt_3041_branch_req_0 : boolean;
  signal SUB_u32_u32_3071_inst_req_0 : boolean;
  signal ADD_u32_u32_3104_inst_ack_1 : boolean;
  signal ULT_u32_u1_2876_inst_req_0 : boolean;
  signal ULT_u32_u1_2876_inst_ack_0 : boolean;
  signal ULT_u32_u1_2876_inst_req_1 : boolean;
  signal ULT_u32_u1_2876_inst_ack_1 : boolean;
  signal ADD_u32_u32_3104_inst_req_1 : boolean;
  signal OR_u32_u32_3114_inst_ack_0 : boolean;
  signal if_stmt_2878_branch_req_0 : boolean;
  signal if_stmt_2878_branch_ack_1 : boolean;
  signal if_stmt_2878_branch_ack_0 : boolean;
  signal AND_u32_u32_3092_inst_ack_1 : boolean;
  signal SUB_u32_u32_3066_inst_ack_0 : boolean;
  signal SUB_u32_u32_3071_inst_req_1 : boolean;
  signal SUB_u32_u32_3066_inst_req_1 : boolean;
  signal ADD_u32_u32_3039_inst_ack_1 : boolean;
  signal ADD_u32_u32_3061_inst_ack_1 : boolean;
  signal ADD_u32_u32_3039_inst_req_1 : boolean;
  signal ADD_u32_u32_2913_inst_req_0 : boolean;
  signal ADD_u32_u32_2913_inst_ack_0 : boolean;
  signal ADD_u32_u32_2913_inst_req_1 : boolean;
  signal ADD_u32_u32_2913_inst_ack_1 : boolean;
  signal OR_u32_u32_3114_inst_req_0 : boolean;
  signal SUB_u32_u32_3066_inst_req_0 : boolean;
  signal AND_u32_u32_3092_inst_req_0 : boolean;
  signal ADD_u32_u32_3039_inst_ack_0 : boolean;
  signal SUB_u32_u32_2918_inst_req_0 : boolean;
  signal SUB_u32_u32_2918_inst_ack_0 : boolean;
  signal ADD_u32_u32_3039_inst_req_0 : boolean;
  signal SUB_u32_u32_2918_inst_req_1 : boolean;
  signal SUB_u32_u32_2918_inst_ack_1 : boolean;
  signal ADD_u32_u32_3104_inst_ack_0 : boolean;
  signal ADD_u32_u32_3104_inst_req_0 : boolean;
  signal ULT_u32_u1_2923_inst_req_0 : boolean;
  signal ULT_u32_u1_2923_inst_ack_0 : boolean;
  signal ULT_u32_u1_2923_inst_req_1 : boolean;
  signal ULT_u32_u1_2923_inst_ack_1 : boolean;
  signal if_stmt_2925_branch_req_0 : boolean;
  signal if_stmt_2925_branch_ack_1 : boolean;
  signal if_stmt_2925_branch_ack_0 : boolean;
  signal type_cast_3024_inst_req_1 : boolean;
  signal AND_u32_u32_2960_inst_req_0 : boolean;
  signal AND_u32_u32_2960_inst_ack_0 : boolean;
  signal AND_u1_u1_3033_inst_ack_1 : boolean;
  signal AND_u32_u32_2960_inst_req_1 : boolean;
  signal AND_u32_u32_2960_inst_ack_1 : boolean;
  signal AND_u1_u1_3033_inst_req_1 : boolean;
  signal ADD_u32_u32_3061_inst_req_0 : boolean;
  signal SHL_u32_u32_3098_inst_ack_1 : boolean;
  signal AND_u1_u1_3033_inst_ack_0 : boolean;
  signal EQ_u32_u1_2966_inst_req_0 : boolean;
  signal EQ_u32_u1_2966_inst_ack_0 : boolean;
  signal AND_u1_u1_3033_inst_req_0 : boolean;
  signal EQ_u32_u1_2966_inst_req_1 : boolean;
  signal EQ_u32_u1_2966_inst_ack_1 : boolean;
  signal SHL_u32_u32_3098_inst_req_1 : boolean;
  signal ADD_u32_u32_3061_inst_req_1 : boolean;
  signal type_cast_2970_inst_req_0 : boolean;
  signal type_cast_2970_inst_ack_0 : boolean;
  signal type_cast_2970_inst_req_1 : boolean;
  signal type_cast_2970_inst_ack_1 : boolean;
  signal SUB_u32_u32_3071_inst_ack_1 : boolean;
  signal NEQ_i32_u1_2974_inst_req_0 : boolean;
  signal NEQ_i32_u1_2974_inst_ack_0 : boolean;
  signal NEQ_i32_u1_2974_inst_req_1 : boolean;
  signal NEQ_i32_u1_2974_inst_ack_1 : boolean;
  signal SUB_u32_u32_3066_inst_ack_1 : boolean;
  signal AND_u1_u1_2979_inst_req_0 : boolean;
  signal AND_u1_u1_2979_inst_ack_0 : boolean;
  signal AND_u1_u1_2979_inst_req_1 : boolean;
  signal AND_u1_u1_2979_inst_ack_1 : boolean;
  signal OR_u32_u32_3109_inst_ack_1 : boolean;
  signal EQ_u32_u1_3020_inst_ack_1 : boolean;
  signal NEQ_i32_u1_3028_inst_ack_1 : boolean;
  signal if_stmt_2981_branch_req_0 : boolean;
  signal if_stmt_2981_branch_ack_1 : boolean;
  signal if_stmt_2981_branch_ack_0 : boolean;
  signal SHL_u32_u32_3008_inst_req_0 : boolean;
  signal SHL_u32_u32_3008_inst_ack_0 : boolean;
  signal SHL_u32_u32_3008_inst_req_1 : boolean;
  signal SHL_u32_u32_3008_inst_ack_1 : boolean;
  signal AND_u32_u32_3014_inst_req_0 : boolean;
  signal AND_u32_u32_3014_inst_ack_0 : boolean;
  signal AND_u32_u32_3014_inst_req_1 : boolean;
  signal AND_u32_u32_3014_inst_ack_1 : boolean;
  signal EQ_u32_u1_3020_inst_req_0 : boolean;
  signal EQ_u32_u1_3020_inst_ack_0 : boolean;
  signal EQ_u32_u1_3020_inst_req_1 : boolean;
  signal type_cast_3118_inst_req_0 : boolean;
  signal type_cast_3118_inst_ack_0 : boolean;
  signal type_cast_3118_inst_req_1 : boolean;
  signal type_cast_3118_inst_ack_1 : boolean;
  signal SLT_f32_u1_3134_inst_req_0 : boolean;
  signal SLT_f32_u1_3134_inst_ack_0 : boolean;
  signal SLT_f32_u1_3134_inst_req_1 : boolean;
  signal SLT_f32_u1_3134_inst_ack_1 : boolean;
  signal MUL_f32_f32_3140_inst_req_0 : boolean;
  signal MUL_f32_f32_3140_inst_ack_0 : boolean;
  signal MUL_f32_f32_3140_inst_req_1 : boolean;
  signal MUL_f32_f32_3140_inst_ack_1 : boolean;
  signal type_cast_3144_inst_req_0 : boolean;
  signal type_cast_3144_inst_ack_0 : boolean;
  signal type_cast_3144_inst_req_1 : boolean;
  signal type_cast_3144_inst_ack_1 : boolean;
  signal type_cast_3148_inst_req_0 : boolean;
  signal type_cast_3148_inst_ack_0 : boolean;
  signal type_cast_3148_inst_req_1 : boolean;
  signal type_cast_3148_inst_ack_1 : boolean;
  signal MUX_3155_inst_req_0 : boolean;
  signal MUX_3155_inst_ack_0 : boolean;
  signal MUX_3155_inst_req_1 : boolean;
  signal MUX_3155_inst_ack_1 : boolean;
  signal EQ_f32_u1_3161_inst_req_0 : boolean;
  signal EQ_f32_u1_3161_inst_ack_0 : boolean;
  signal EQ_f32_u1_3161_inst_req_1 : boolean;
  signal EQ_f32_u1_3161_inst_ack_1 : boolean;
  signal if_stmt_3163_branch_req_0 : boolean;
  signal if_stmt_3163_branch_ack_1 : boolean;
  signal if_stmt_3163_branch_ack_0 : boolean;
  signal LSHR_u32_u32_3174_inst_req_0 : boolean;
  signal LSHR_u32_u32_3174_inst_ack_0 : boolean;
  signal LSHR_u32_u32_3174_inst_req_1 : boolean;
  signal LSHR_u32_u32_3174_inst_ack_1 : boolean;
  signal AND_u32_u32_3180_inst_req_0 : boolean;
  signal AND_u32_u32_3180_inst_ack_0 : boolean;
  signal AND_u32_u32_3180_inst_req_1 : boolean;
  signal AND_u32_u32_3180_inst_ack_1 : boolean;
  signal LSHR_u32_u32_3186_inst_req_0 : boolean;
  signal LSHR_u32_u32_3186_inst_ack_0 : boolean;
  signal LSHR_u32_u32_3186_inst_req_1 : boolean;
  signal LSHR_u32_u32_3186_inst_ack_1 : boolean;
  signal AND_u32_u32_3192_inst_req_0 : boolean;
  signal AND_u32_u32_3192_inst_ack_0 : boolean;
  signal AND_u32_u32_3192_inst_req_1 : boolean;
  signal AND_u32_u32_3192_inst_ack_1 : boolean;
  signal if_stmt_3838_branch_ack_1 : boolean;
  signal SHL_u32_u32_3198_inst_req_0 : boolean;
  signal SHL_u32_u32_3198_inst_ack_0 : boolean;
  signal SHL_u32_u32_3198_inst_req_1 : boolean;
  signal SHL_u32_u32_3198_inst_ack_1 : boolean;
  signal if_stmt_3789_branch_ack_0 : boolean;
  signal ADD_u32_u32_3825_inst_req_0 : boolean;
  signal AND_u32_u32_3204_inst_req_0 : boolean;
  signal AND_u32_u32_3204_inst_ack_0 : boolean;
  signal AND_u32_u32_3204_inst_req_1 : boolean;
  signal AND_u32_u32_3204_inst_ack_1 : boolean;
  signal ADD_u32_u32_3825_inst_ack_0 : boolean;
  signal OR_u32_u32_3210_inst_req_0 : boolean;
  signal OR_u32_u32_3210_inst_ack_0 : boolean;
  signal OR_u32_u32_3210_inst_req_1 : boolean;
  signal OR_u32_u32_3210_inst_ack_1 : boolean;
  signal LSHR_u32_u32_3216_inst_req_0 : boolean;
  signal LSHR_u32_u32_3216_inst_ack_0 : boolean;
  signal LSHR_u32_u32_3216_inst_req_1 : boolean;
  signal LSHR_u32_u32_3216_inst_ack_1 : boolean;
  signal AND_u32_u32_3222_inst_req_0 : boolean;
  signal AND_u32_u32_3222_inst_ack_0 : boolean;
  signal AND_u32_u32_3222_inst_req_1 : boolean;
  signal AND_u32_u32_3222_inst_ack_1 : boolean;
  signal if_stmt_3789_branch_ack_1 : boolean;
  signal OR_u32_u32_3228_inst_req_0 : boolean;
  signal OR_u32_u32_3228_inst_ack_0 : boolean;
  signal OR_u32_u32_3228_inst_req_1 : boolean;
  signal OR_u32_u32_3228_inst_ack_1 : boolean;
  signal ADD_u32_u32_3825_inst_req_1 : boolean;
  signal SUB_u32_u32_3830_inst_req_1 : boolean;
  signal XOR_u32_u32_3233_inst_req_0 : boolean;
  signal XOR_u32_u32_3233_inst_ack_0 : boolean;
  signal XOR_u32_u32_3233_inst_req_1 : boolean;
  signal XOR_u32_u32_3233_inst_ack_1 : boolean;
  signal ADD_u32_u32_3825_inst_ack_1 : boolean;
  signal if_stmt_3838_branch_ack_0 : boolean;
  signal AND_u32_u32_3239_inst_req_0 : boolean;
  signal AND_u32_u32_3239_inst_ack_0 : boolean;
  signal AND_u32_u32_3239_inst_req_1 : boolean;
  signal AND_u32_u32_3239_inst_ack_1 : boolean;
  signal SUB_u32_u32_3244_inst_req_0 : boolean;
  signal SUB_u32_u32_3244_inst_ack_0 : boolean;
  signal SUB_u32_u32_3244_inst_req_1 : boolean;
  signal SUB_u32_u32_3244_inst_ack_1 : boolean;
  signal switch_stmt_3246_branch_default_req_0 : boolean;
  signal switch_stmt_3246_select_expr_0_req_0 : boolean;
  signal switch_stmt_3246_select_expr_0_ack_0 : boolean;
  signal switch_stmt_3246_select_expr_0_req_1 : boolean;
  signal switch_stmt_3246_select_expr_0_ack_1 : boolean;
  signal switch_stmt_3246_branch_0_req_0 : boolean;
  signal switch_stmt_3246_select_expr_1_req_0 : boolean;
  signal switch_stmt_3246_select_expr_1_ack_0 : boolean;
  signal switch_stmt_3246_select_expr_1_req_1 : boolean;
  signal switch_stmt_3246_select_expr_1_ack_1 : boolean;
  signal switch_stmt_3246_branch_1_req_0 : boolean;
  signal switch_stmt_3246_branch_0_ack_1 : boolean;
  signal switch_stmt_3246_branch_1_ack_1 : boolean;
  signal SUB_u32_u32_3830_inst_req_0 : boolean;
  signal switch_stmt_3246_branch_default_ack_0 : boolean;
  signal SUB_u32_u32_3830_inst_ack_0 : boolean;
  signal ULT_u32_u1_3836_inst_req_1 : boolean;
  signal LSHR_u32_u32_3277_inst_req_0 : boolean;
  signal LSHR_u32_u32_3277_inst_ack_0 : boolean;
  signal LSHR_u32_u32_3277_inst_req_1 : boolean;
  signal LSHR_u32_u32_3277_inst_ack_1 : boolean;
  signal if_stmt_3838_branch_req_0 : boolean;
  signal ULT_u32_u1_3836_inst_req_0 : boolean;
  signal ULT_u32_u1_3836_inst_ack_1 : boolean;
  signal UGT_u32_u1_3282_inst_req_0 : boolean;
  signal UGT_u32_u1_3282_inst_ack_0 : boolean;
  signal UGT_u32_u1_3282_inst_req_1 : boolean;
  signal UGT_u32_u1_3282_inst_ack_1 : boolean;
  signal ULT_u32_u1_3836_inst_ack_0 : boolean;
  signal if_stmt_3284_branch_req_0 : boolean;
  signal if_stmt_3284_branch_ack_1 : boolean;
  signal if_stmt_3284_branch_ack_0 : boolean;
  signal if_stmt_3789_branch_req_0 : boolean;
  signal SHL_u32_u32_3311_inst_req_0 : boolean;
  signal SHL_u32_u32_3311_inst_ack_0 : boolean;
  signal SHL_u32_u32_3311_inst_req_1 : boolean;
  signal SHL_u32_u32_3311_inst_ack_1 : boolean;
  signal SUB_u32_u32_3830_inst_ack_1 : boolean;
  signal SHL_u32_u32_3317_inst_req_0 : boolean;
  signal SHL_u32_u32_3317_inst_ack_0 : boolean;
  signal SHL_u32_u32_3317_inst_req_1 : boolean;
  signal SHL_u32_u32_3317_inst_ack_1 : boolean;
  signal ULT_u32_u1_3322_inst_req_0 : boolean;
  signal ULT_u32_u1_3322_inst_ack_0 : boolean;
  signal ULT_u32_u1_3322_inst_req_1 : boolean;
  signal ULT_u32_u1_3322_inst_ack_1 : boolean;
  signal if_stmt_3324_branch_req_0 : boolean;
  signal if_stmt_3324_branch_ack_1 : boolean;
  signal if_stmt_3324_branch_ack_0 : boolean;
  signal ADD_u32_u32_3359_inst_req_0 : boolean;
  signal ADD_u32_u32_3359_inst_ack_0 : boolean;
  signal ADD_u32_u32_3359_inst_req_1 : boolean;
  signal ADD_u32_u32_3359_inst_ack_1 : boolean;
  signal SUB_u32_u32_3364_inst_req_0 : boolean;
  signal SUB_u32_u32_3364_inst_ack_0 : boolean;
  signal SUB_u32_u32_3364_inst_req_1 : boolean;
  signal SUB_u32_u32_3364_inst_ack_1 : boolean;
  signal ULT_u32_u1_3369_inst_req_0 : boolean;
  signal ULT_u32_u1_3369_inst_ack_0 : boolean;
  signal ULT_u32_u1_3369_inst_req_1 : boolean;
  signal ULT_u32_u1_3369_inst_ack_1 : boolean;
  signal if_stmt_3371_branch_req_0 : boolean;
  signal if_stmt_3371_branch_ack_1 : boolean;
  signal if_stmt_3371_branch_ack_0 : boolean;
  signal AND_u32_u32_3406_inst_req_0 : boolean;
  signal AND_u32_u32_3406_inst_ack_0 : boolean;
  signal AND_u32_u32_3406_inst_req_1 : boolean;
  signal AND_u32_u32_3406_inst_ack_1 : boolean;
  signal EQ_u32_u1_3412_inst_req_0 : boolean;
  signal EQ_u32_u1_3412_inst_ack_0 : boolean;
  signal EQ_u32_u1_3412_inst_req_1 : boolean;
  signal EQ_u32_u1_3412_inst_ack_1 : boolean;
  signal type_cast_3416_inst_req_0 : boolean;
  signal type_cast_3416_inst_ack_0 : boolean;
  signal type_cast_3416_inst_req_1 : boolean;
  signal type_cast_3416_inst_ack_1 : boolean;
  signal NEQ_i32_u1_3420_inst_req_0 : boolean;
  signal NEQ_i32_u1_3420_inst_ack_0 : boolean;
  signal NEQ_i32_u1_3420_inst_req_1 : boolean;
  signal NEQ_i32_u1_3420_inst_ack_1 : boolean;
  signal AND_u1_u1_3425_inst_req_0 : boolean;
  signal AND_u1_u1_3425_inst_ack_0 : boolean;
  signal AND_u1_u1_3425_inst_req_1 : boolean;
  signal AND_u1_u1_3425_inst_ack_1 : boolean;
  signal if_stmt_3427_branch_req_0 : boolean;
  signal if_stmt_3427_branch_ack_1 : boolean;
  signal if_stmt_3427_branch_ack_0 : boolean;
  signal SHL_u32_u32_3454_inst_req_0 : boolean;
  signal SHL_u32_u32_3454_inst_ack_0 : boolean;
  signal SHL_u32_u32_3454_inst_req_1 : boolean;
  signal SHL_u32_u32_3454_inst_ack_1 : boolean;
  signal AND_u32_u32_3460_inst_req_0 : boolean;
  signal EQ_u32_u1_3466_inst_req_0 : boolean;
  signal EQ_u32_u1_3466_inst_ack_0 : boolean;
  signal EQ_u32_u1_3466_inst_req_1 : boolean;
  signal EQ_u32_u1_3466_inst_ack_1 : boolean;
  signal type_cast_3470_inst_req_0 : boolean;
  signal type_cast_3470_inst_ack_0 : boolean;
  signal type_cast_3470_inst_req_1 : boolean;
  signal type_cast_3470_inst_ack_1 : boolean;
  signal NEQ_i32_u1_3474_inst_req_0 : boolean;
  signal NEQ_i32_u1_3474_inst_ack_0 : boolean;
  signal NEQ_i32_u1_3474_inst_req_1 : boolean;
  signal NEQ_i32_u1_3474_inst_ack_1 : boolean;
  signal AND_u1_u1_3479_inst_req_0 : boolean;
  signal AND_u1_u1_3479_inst_ack_0 : boolean;
  signal AND_u1_u1_3479_inst_req_1 : boolean;
  signal AND_u1_u1_3479_inst_ack_1 : boolean;
  signal ADD_u32_u32_3485_inst_req_0 : boolean;
  signal ADD_u32_u32_3485_inst_ack_0 : boolean;
  signal ADD_u32_u32_3485_inst_req_1 : boolean;
  signal ADD_u32_u32_3485_inst_ack_1 : boolean;
  signal if_stmt_3487_branch_req_0 : boolean;
  signal if_stmt_3487_branch_ack_1 : boolean;
  signal if_stmt_3487_branch_ack_0 : boolean;
  signal ADD_u32_u32_3507_inst_req_0 : boolean;
  signal ADD_u32_u32_3507_inst_ack_0 : boolean;
  signal ADD_u32_u32_3507_inst_req_1 : boolean;
  signal ADD_u32_u32_3507_inst_ack_1 : boolean;
  signal SUB_u32_u32_3512_inst_req_0 : boolean;
  signal SUB_u32_u32_3512_inst_ack_0 : boolean;
  signal SUB_u32_u32_3512_inst_req_1 : boolean;
  signal SUB_u32_u32_3512_inst_ack_1 : boolean;
  signal SUB_u32_u32_3517_inst_req_0 : boolean;
  signal SUB_u32_u32_3517_inst_ack_0 : boolean;
  signal SUB_u32_u32_3517_inst_req_1 : boolean;
  signal SUB_u32_u32_3517_inst_ack_1 : boolean;
  signal AND_u32_u32_3538_inst_req_0 : boolean;
  signal AND_u32_u32_3538_inst_ack_0 : boolean;
  signal AND_u32_u32_3538_inst_req_1 : boolean;
  signal AND_u32_u32_3538_inst_ack_1 : boolean;
  signal SHL_u32_u32_3544_inst_req_0 : boolean;
  signal SHL_u32_u32_3544_inst_ack_0 : boolean;
  signal SHL_u32_u32_3544_inst_req_1 : boolean;
  signal SHL_u32_u32_3544_inst_ack_1 : boolean;
  signal ADD_u32_u32_3550_inst_req_0 : boolean;
  signal ADD_u32_u32_3550_inst_ack_0 : boolean;
  signal ADD_u32_u32_3550_inst_req_1 : boolean;
  signal ADD_u32_u32_3550_inst_ack_1 : boolean;
  signal OR_u32_u32_3555_inst_req_0 : boolean;
  signal OR_u32_u32_3555_inst_ack_0 : boolean;
  signal OR_u32_u32_3555_inst_req_1 : boolean;
  signal OR_u32_u32_3555_inst_ack_1 : boolean;
  signal OR_u32_u32_3560_inst_req_0 : boolean;
  signal OR_u32_u32_3560_inst_ack_0 : boolean;
  signal OR_u32_u32_3560_inst_req_1 : boolean;
  signal OR_u32_u32_3560_inst_ack_1 : boolean;
  signal type_cast_3564_inst_req_0 : boolean;
  signal type_cast_3564_inst_ack_0 : boolean;
  signal type_cast_3564_inst_req_1 : boolean;
  signal type_cast_3564_inst_ack_1 : boolean;
  signal SUB_f32_f32_3579_inst_req_0 : boolean;
  signal SUB_f32_f32_3579_inst_ack_0 : boolean;
  signal SUB_f32_f32_3579_inst_req_1 : boolean;
  signal SUB_f32_f32_3579_inst_ack_1 : boolean;
  signal WPIPE_out_data_4043_inst_ack_0 : boolean;
  signal MUL_f32_f32_3585_inst_req_0 : boolean;
  signal MUL_f32_f32_3585_inst_ack_0 : boolean;
  signal MUL_f32_f32_3585_inst_req_1 : boolean;
  signal MUL_f32_f32_3585_inst_ack_1 : boolean;
  signal WPIPE_out_data_4052_inst_ack_1 : boolean;
  signal ADD_f32_f32_3590_inst_req_0 : boolean;
  signal ADD_f32_f32_3590_inst_ack_0 : boolean;
  signal ADD_f32_f32_3590_inst_req_1 : boolean;
  signal ADD_f32_f32_3590_inst_ack_1 : boolean;
  signal WPIPE_out_data_4043_inst_req_1 : boolean;
  signal phi_stmt_2045_req_0 : boolean;
  signal MUL_f32_f32_3596_inst_req_0 : boolean;
  signal MUL_f32_f32_3596_inst_ack_0 : boolean;
  signal MUL_f32_f32_3596_inst_req_1 : boolean;
  signal MUL_f32_f32_3596_inst_ack_1 : boolean;
  signal SLT_f32_u1_3602_inst_req_0 : boolean;
  signal SLT_f32_u1_3602_inst_ack_0 : boolean;
  signal SLT_f32_u1_3602_inst_req_1 : boolean;
  signal SLT_f32_u1_3602_inst_ack_1 : boolean;
  signal WPIPE_out_data_4043_inst_ack_1 : boolean;
  signal if_stmt_3604_branch_req_0 : boolean;
  signal type_cast_4031_inst_req_1 : boolean;
  signal if_stmt_3604_branch_ack_1 : boolean;
  signal if_stmt_3604_branch_ack_0 : boolean;
  signal type_cast_4031_inst_ack_1 : boolean;
  signal phi_stmt_2052_req_0 : boolean;
  signal SGT_f32_u1_3615_inst_req_0 : boolean;
  signal SGT_f32_u1_3615_inst_ack_0 : boolean;
  signal SGT_f32_u1_3615_inst_req_1 : boolean;
  signal SGT_f32_u1_3615_inst_ack_1 : boolean;
  signal if_stmt_3617_branch_req_0 : boolean;
  signal if_stmt_3617_branch_ack_1 : boolean;
  signal if_stmt_3617_branch_ack_0 : boolean;
  signal MUL_f32_f32_3641_inst_req_0 : boolean;
  signal MUL_f32_f32_3641_inst_ack_0 : boolean;
  signal MUL_f32_f32_3641_inst_req_1 : boolean;
  signal MUL_f32_f32_3641_inst_ack_1 : boolean;
  signal type_cast_2065_inst_req_0 : boolean;
  signal type_cast_2065_inst_ack_0 : boolean;
  signal ADD_f32_f32_3646_inst_req_0 : boolean;
  signal ADD_f32_f32_3646_inst_ack_0 : boolean;
  signal ADD_f32_f32_3646_inst_req_1 : boolean;
  signal ADD_f32_f32_3646_inst_ack_1 : boolean;
  signal SLT_f32_u1_3652_inst_req_0 : boolean;
  signal SLT_f32_u1_3652_inst_ack_0 : boolean;
  signal SLT_f32_u1_3652_inst_req_1 : boolean;
  signal SLT_f32_u1_3652_inst_ack_1 : boolean;
  signal if_stmt_3654_branch_req_0 : boolean;
  signal if_stmt_3654_branch_ack_1 : boolean;
  signal if_stmt_3654_branch_ack_0 : boolean;
  signal SGT_f32_u1_3665_inst_req_0 : boolean;
  signal SGT_f32_u1_3665_inst_ack_0 : boolean;
  signal SGT_f32_u1_3665_inst_req_1 : boolean;
  signal SGT_f32_u1_3665_inst_ack_1 : boolean;
  signal if_stmt_3667_branch_req_0 : boolean;
  signal if_stmt_3667_branch_ack_1 : boolean;
  signal if_stmt_3667_branch_ack_0 : boolean;
  signal EQ_f32_u1_3678_inst_req_0 : boolean;
  signal EQ_f32_u1_3678_inst_ack_0 : boolean;
  signal EQ_f32_u1_3678_inst_req_1 : boolean;
  signal EQ_f32_u1_3678_inst_ack_1 : boolean;
  signal if_stmt_3680_branch_req_0 : boolean;
  signal if_stmt_3680_branch_ack_1 : boolean;
  signal if_stmt_3680_branch_ack_0 : boolean;
  signal type_cast_3700_inst_req_0 : boolean;
  signal type_cast_3700_inst_ack_0 : boolean;
  signal type_cast_3700_inst_req_1 : boolean;
  signal type_cast_3700_inst_ack_1 : boolean;
  signal SHL_u32_u32_3706_inst_req_0 : boolean;
  signal SHL_u32_u32_3706_inst_ack_0 : boolean;
  signal SHL_u32_u32_3706_inst_req_1 : boolean;
  signal SHL_u32_u32_3706_inst_ack_1 : boolean;
  signal AND_u32_u32_3712_inst_req_0 : boolean;
  signal AND_u32_u32_3712_inst_ack_0 : boolean;
  signal AND_u32_u32_3712_inst_req_1 : boolean;
  signal AND_u32_u32_3712_inst_ack_1 : boolean;
  signal OR_u32_u32_3718_inst_req_0 : boolean;
  signal OR_u32_u32_3718_inst_ack_0 : boolean;
  signal OR_u32_u32_3718_inst_req_1 : boolean;
  signal OR_u32_u32_3718_inst_ack_1 : boolean;
  signal LSHR_u32_u32_3740_inst_req_0 : boolean;
  signal LSHR_u32_u32_3740_inst_ack_0 : boolean;
  signal LSHR_u32_u32_3740_inst_req_1 : boolean;
  signal LSHR_u32_u32_3740_inst_ack_1 : boolean;
  signal UGT_u32_u1_3746_inst_req_0 : boolean;
  signal UGT_u32_u1_3746_inst_ack_0 : boolean;
  signal UGT_u32_u1_3746_inst_req_1 : boolean;
  signal UGT_u32_u1_3746_inst_ack_1 : boolean;
  signal if_stmt_3748_branch_req_0 : boolean;
  signal if_stmt_3748_branch_ack_1 : boolean;
  signal if_stmt_3748_branch_ack_0 : boolean;
  signal SHL_u32_u32_3776_inst_req_0 : boolean;
  signal SHL_u32_u32_3776_inst_ack_0 : boolean;
  signal SHL_u32_u32_3776_inst_req_1 : boolean;
  signal SHL_u32_u32_3776_inst_ack_1 : boolean;
  signal SHL_u32_u32_3782_inst_req_0 : boolean;
  signal SHL_u32_u32_3782_inst_ack_0 : boolean;
  signal SHL_u32_u32_3782_inst_req_1 : boolean;
  signal SHL_u32_u32_3782_inst_ack_1 : boolean;
  signal ULT_u32_u1_3787_inst_req_0 : boolean;
  signal ULT_u32_u1_3787_inst_ack_0 : boolean;
  signal ULT_u32_u1_3787_inst_req_1 : boolean;
  signal ULT_u32_u1_3787_inst_ack_1 : boolean;
  signal LSHR_u32_u32_3854_inst_req_0 : boolean;
  signal LSHR_u32_u32_3854_inst_ack_0 : boolean;
  signal LSHR_u32_u32_3854_inst_req_1 : boolean;
  signal LSHR_u32_u32_3854_inst_ack_1 : boolean;
  signal AND_u32_u32_3860_inst_req_0 : boolean;
  signal AND_u32_u32_3860_inst_ack_0 : boolean;
  signal AND_u32_u32_3860_inst_req_1 : boolean;
  signal AND_u32_u32_3860_inst_ack_1 : boolean;
  signal AND_u32_u32_3866_inst_req_0 : boolean;
  signal AND_u32_u32_3866_inst_ack_0 : boolean;
  signal AND_u32_u32_3866_inst_req_1 : boolean;
  signal AND_u32_u32_3866_inst_ack_1 : boolean;
  signal ADD_u32_u32_3872_inst_req_0 : boolean;
  signal ADD_u32_u32_3872_inst_ack_0 : boolean;
  signal ADD_u32_u32_3872_inst_req_1 : boolean;
  signal ADD_u32_u32_3872_inst_ack_1 : boolean;
  signal AND_u32_u32_3878_inst_req_0 : boolean;
  signal AND_u32_u32_3878_inst_ack_0 : boolean;
  signal AND_u32_u32_3878_inst_req_1 : boolean;
  signal AND_u32_u32_3878_inst_ack_1 : boolean;
  signal EQ_u32_u1_3884_inst_req_0 : boolean;
  signal EQ_u32_u1_3884_inst_ack_0 : boolean;
  signal EQ_u32_u1_3884_inst_req_1 : boolean;
  signal EQ_u32_u1_3884_inst_ack_1 : boolean;
  signal type_cast_3888_inst_req_0 : boolean;
  signal type_cast_3888_inst_ack_0 : boolean;
  signal type_cast_3888_inst_req_1 : boolean;
  signal type_cast_3888_inst_ack_1 : boolean;
  signal NEQ_i32_u1_3892_inst_req_0 : boolean;
  signal NEQ_i32_u1_3892_inst_ack_0 : boolean;
  signal NEQ_i32_u1_3892_inst_req_1 : boolean;
  signal NEQ_i32_u1_3892_inst_ack_1 : boolean;
  signal AND_u1_u1_3897_inst_req_0 : boolean;
  signal AND_u1_u1_3897_inst_ack_0 : boolean;
  signal AND_u1_u1_3897_inst_req_1 : boolean;
  signal AND_u1_u1_3897_inst_ack_1 : boolean;
  signal if_stmt_3899_branch_req_0 : boolean;
  signal if_stmt_3899_branch_ack_1 : boolean;
  signal if_stmt_3899_branch_ack_0 : boolean;
  signal SHL_u32_u32_3926_inst_req_0 : boolean;
  signal SHL_u32_u32_3926_inst_ack_0 : boolean;
  signal SHL_u32_u32_3926_inst_req_1 : boolean;
  signal SHL_u32_u32_3926_inst_ack_1 : boolean;
  signal AND_u32_u32_3932_inst_req_0 : boolean;
  signal AND_u32_u32_3932_inst_ack_0 : boolean;
  signal AND_u32_u32_3932_inst_req_1 : boolean;
  signal AND_u32_u32_3932_inst_ack_1 : boolean;
  signal WPIPE_out_data_4052_inst_req_1 : boolean;
  signal WPIPE_out_data_4052_inst_ack_0 : boolean;
  signal EQ_u32_u1_3938_inst_req_0 : boolean;
  signal EQ_u32_u1_3938_inst_ack_0 : boolean;
  signal WPIPE_out_data_4052_inst_req_0 : boolean;
  signal EQ_u32_u1_3938_inst_req_1 : boolean;
  signal EQ_u32_u1_3938_inst_ack_1 : boolean;
  signal phi_stmt_2045_req_1 : boolean;
  signal phi_stmt_2059_ack_0 : boolean;
  signal type_cast_2051_inst_ack_1 : boolean;
  signal type_cast_2051_inst_req_1 : boolean;
  signal type_cast_3942_inst_req_0 : boolean;
  signal type_cast_3942_inst_ack_0 : boolean;
  signal type_cast_3942_inst_req_1 : boolean;
  signal type_cast_3942_inst_ack_1 : boolean;
  signal phi_stmt_2045_ack_0 : boolean;
  signal phi_stmt_2052_ack_0 : boolean;
  signal type_cast_2051_inst_ack_0 : boolean;
  signal type_cast_2051_inst_req_0 : boolean;
  signal NEQ_i32_u1_3946_inst_req_0 : boolean;
  signal NEQ_i32_u1_3946_inst_ack_0 : boolean;
  signal NEQ_i32_u1_3946_inst_req_1 : boolean;
  signal NEQ_i32_u1_3946_inst_ack_1 : boolean;
  signal phi_stmt_2059_req_0 : boolean;
  signal WPIPE_out_data_4049_inst_ack_1 : boolean;
  signal WPIPE_out_data_4049_inst_req_1 : boolean;
  signal AND_u1_u1_3951_inst_req_0 : boolean;
  signal AND_u1_u1_3951_inst_ack_0 : boolean;
  signal AND_u1_u1_3951_inst_req_1 : boolean;
  signal AND_u1_u1_3951_inst_ack_1 : boolean;
  signal phi_stmt_2059_req_1 : boolean;
  signal WPIPE_out_data_4049_inst_ack_0 : boolean;
  signal WPIPE_out_data_4043_inst_req_0 : boolean;
  signal WPIPE_out_data_4049_inst_req_0 : boolean;
  signal ADD_u32_u32_3957_inst_req_0 : boolean;
  signal ADD_u32_u32_3957_inst_ack_0 : boolean;
  signal ADD_u32_u32_3957_inst_req_1 : boolean;
  signal ADD_u32_u32_3957_inst_ack_1 : boolean;
  signal phi_stmt_2052_req_1 : boolean;
  signal type_cast_4031_inst_ack_0 : boolean;
  signal if_stmt_3959_branch_req_0 : boolean;
  signal type_cast_4031_inst_req_0 : boolean;
  signal if_stmt_3959_branch_ack_1 : boolean;
  signal if_stmt_3959_branch_ack_0 : boolean;
  signal type_cast_2065_inst_req_1 : boolean;
  signal type_cast_2065_inst_ack_1 : boolean;
  signal type_cast_2058_inst_ack_1 : boolean;
  signal type_cast_2058_inst_req_1 : boolean;
  signal ADD_u32_u32_3979_inst_req_0 : boolean;
  signal ADD_u32_u32_3979_inst_ack_0 : boolean;
  signal ADD_u32_u32_3979_inst_req_1 : boolean;
  signal ADD_u32_u32_3979_inst_ack_1 : boolean;
  signal type_cast_2058_inst_ack_0 : boolean;
  signal type_cast_2058_inst_req_0 : boolean;
  signal WPIPE_out_data_4046_inst_ack_1 : boolean;
  signal SUB_u32_u32_3984_inst_req_0 : boolean;
  signal SUB_u32_u32_3984_inst_ack_0 : boolean;
  signal WPIPE_out_data_4046_inst_req_1 : boolean;
  signal SUB_u32_u32_3984_inst_req_1 : boolean;
  signal SUB_u32_u32_3984_inst_ack_1 : boolean;
  signal AND_u32_u32_4005_inst_req_0 : boolean;
  signal AND_u32_u32_4005_inst_ack_0 : boolean;
  signal WPIPE_out_data_4046_inst_ack_0 : boolean;
  signal AND_u32_u32_4005_inst_req_1 : boolean;
  signal AND_u32_u32_4005_inst_ack_1 : boolean;
  signal WPIPE_out_data_4046_inst_req_0 : boolean;
  signal SHL_u32_u32_4011_inst_req_0 : boolean;
  signal SHL_u32_u32_4011_inst_ack_0 : boolean;
  signal SHL_u32_u32_4011_inst_req_1 : boolean;
  signal SHL_u32_u32_4011_inst_ack_1 : boolean;
  signal ADD_u32_u32_4017_inst_req_0 : boolean;
  signal ADD_u32_u32_4017_inst_ack_0 : boolean;
  signal ADD_u32_u32_4017_inst_req_1 : boolean;
  signal ADD_u32_u32_4017_inst_ack_1 : boolean;
  signal OR_u32_u32_4022_inst_req_0 : boolean;
  signal OR_u32_u32_4022_inst_ack_0 : boolean;
  signal OR_u32_u32_4022_inst_req_1 : boolean;
  signal OR_u32_u32_4022_inst_ack_1 : boolean;
  signal phi_stmt_2813_ack_0 : boolean;
  signal phi_stmt_2819_ack_0 : boolean;
  signal OR_u32_u32_4027_inst_req_0 : boolean;
  signal OR_u32_u32_4027_inst_ack_0 : boolean;
  signal OR_u32_u32_4027_inst_req_1 : boolean;
  signal OR_u32_u32_4027_inst_ack_1 : boolean;
  signal phi_stmt_2134_req_1 : boolean;
  signal phi_stmt_2134_req_2 : boolean;
  signal type_cast_2137_inst_req_0 : boolean;
  signal type_cast_2137_inst_ack_0 : boolean;
  signal type_cast_2137_inst_req_1 : boolean;
  signal type_cast_2137_inst_ack_1 : boolean;
  signal phi_stmt_2134_req_0 : boolean;
  signal phi_stmt_2134_ack_0 : boolean;
  signal phi_stmt_2190_req_1 : boolean;
  signal phi_stmt_2190_req_2 : boolean;
  signal type_cast_2193_inst_req_0 : boolean;
  signal type_cast_2193_inst_ack_0 : boolean;
  signal type_cast_2193_inst_req_1 : boolean;
  signal type_cast_2193_inst_ack_1 : boolean;
  signal phi_stmt_2190_req_0 : boolean;
  signal phi_stmt_2190_ack_0 : boolean;
  signal type_cast_2309_inst_req_0 : boolean;
  signal type_cast_2309_inst_ack_0 : boolean;
  signal type_cast_2309_inst_req_1 : boolean;
  signal type_cast_2309_inst_ack_1 : boolean;
  signal phi_stmt_2304_req_1 : boolean;
  signal type_cast_2311_inst_req_0 : boolean;
  signal type_cast_2311_inst_ack_0 : boolean;
  signal type_cast_2311_inst_req_1 : boolean;
  signal type_cast_2311_inst_ack_1 : boolean;
  signal phi_stmt_2304_req_2 : boolean;
  signal phi_stmt_2304_req_3 : boolean;
  signal type_cast_2307_inst_req_0 : boolean;
  signal type_cast_2307_inst_ack_0 : boolean;
  signal type_cast_2307_inst_req_1 : boolean;
  signal type_cast_2307_inst_ack_1 : boolean;
  signal phi_stmt_2304_req_0 : boolean;
  signal phi_stmt_2304_ack_0 : boolean;
  signal type_cast_2375_inst_req_0 : boolean;
  signal type_cast_2375_inst_ack_0 : boolean;
  signal type_cast_2375_inst_req_1 : boolean;
  signal type_cast_2375_inst_ack_1 : boolean;
  signal phi_stmt_2370_req_1 : boolean;
  signal phi_stmt_2376_req_1 : boolean;
  signal type_cast_2373_inst_req_0 : boolean;
  signal type_cast_2373_inst_ack_0 : boolean;
  signal type_cast_2373_inst_req_1 : boolean;
  signal type_cast_2373_inst_ack_1 : boolean;
  signal phi_stmt_2370_req_0 : boolean;
  signal type_cast_2379_inst_req_0 : boolean;
  signal type_cast_2379_inst_ack_0 : boolean;
  signal type_cast_2379_inst_req_1 : boolean;
  signal type_cast_2379_inst_ack_1 : boolean;
  signal phi_stmt_2376_req_0 : boolean;
  signal phi_stmt_2370_ack_0 : boolean;
  signal phi_stmt_2376_ack_0 : boolean;
  signal type_cast_2408_inst_req_0 : boolean;
  signal type_cast_2408_inst_ack_0 : boolean;
  signal type_cast_2408_inst_req_1 : boolean;
  signal type_cast_2408_inst_ack_1 : boolean;
  signal phi_stmt_2405_req_0 : boolean;
  signal type_cast_2415_inst_req_0 : boolean;
  signal type_cast_2415_inst_ack_0 : boolean;
  signal type_cast_2415_inst_req_1 : boolean;
  signal type_cast_2415_inst_ack_1 : boolean;
  signal phi_stmt_2412_req_0 : boolean;
  signal phi_stmt_2405_req_1 : boolean;
  signal phi_stmt_2819_req_0 : boolean;
  signal type_cast_2822_inst_ack_1 : boolean;
  signal type_cast_2822_inst_req_1 : boolean;
  signal phi_stmt_2412_req_1 : boolean;
  signal phi_stmt_2405_ack_0 : boolean;
  signal phi_stmt_2412_ack_0 : boolean;
  signal type_cast_2822_inst_ack_0 : boolean;
  signal type_cast_2822_inst_req_0 : boolean;
  signal type_cast_2447_inst_req_0 : boolean;
  signal type_cast_2447_inst_ack_0 : boolean;
  signal type_cast_2447_inst_req_1 : boolean;
  signal type_cast_2447_inst_ack_1 : boolean;
  signal phi_stmt_2444_req_0 : boolean;
  signal phi_stmt_2813_req_0 : boolean;
  signal type_cast_2451_inst_req_0 : boolean;
  signal type_cast_2451_inst_ack_0 : boolean;
  signal type_cast_2451_inst_req_1 : boolean;
  signal type_cast_2451_inst_ack_1 : boolean;
  signal phi_stmt_2448_req_0 : boolean;
  signal phi_stmt_2444_ack_0 : boolean;
  signal phi_stmt_2448_ack_0 : boolean;
  signal phi_stmt_2455_req_0 : boolean;
  signal type_cast_2816_inst_ack_1 : boolean;
  signal type_cast_2816_inst_req_1 : boolean;
  signal phi_stmt_2462_req_0 : boolean;
  signal type_cast_2816_inst_ack_0 : boolean;
  signal type_cast_2816_inst_req_0 : boolean;
  signal type_cast_2461_inst_req_0 : boolean;
  signal type_cast_2461_inst_ack_0 : boolean;
  signal type_cast_2461_inst_req_1 : boolean;
  signal type_cast_2461_inst_ack_1 : boolean;
  signal phi_stmt_2455_req_1 : boolean;
  signal type_cast_2468_inst_req_0 : boolean;
  signal type_cast_2468_inst_ack_0 : boolean;
  signal type_cast_2468_inst_req_1 : boolean;
  signal type_cast_2468_inst_ack_1 : boolean;
  signal phi_stmt_2462_req_1 : boolean;
  signal phi_stmt_2455_ack_0 : boolean;
  signal phi_stmt_2462_ack_0 : boolean;
  signal phi_stmt_2683_ack_0 : boolean;
  signal type_cast_2496_inst_req_0 : boolean;
  signal type_cast_2496_inst_ack_0 : boolean;
  signal phi_stmt_2819_req_1 : boolean;
  signal type_cast_2496_inst_req_1 : boolean;
  signal type_cast_2496_inst_ack_1 : boolean;
  signal phi_stmt_2493_req_0 : boolean;
  signal phi_stmt_2493_ack_0 : boolean;
  signal phi_stmt_2683_req_0 : boolean;
  signal type_cast_2686_inst_ack_1 : boolean;
  signal type_cast_2559_inst_req_0 : boolean;
  signal type_cast_2559_inst_ack_0 : boolean;
  signal type_cast_2559_inst_req_1 : boolean;
  signal type_cast_2559_inst_ack_1 : boolean;
  signal type_cast_2686_inst_req_1 : boolean;
  signal phi_stmt_2556_req_0 : boolean;
  signal type_cast_2566_inst_req_0 : boolean;
  signal type_cast_2566_inst_ack_0 : boolean;
  signal type_cast_2566_inst_req_1 : boolean;
  signal type_cast_2566_inst_ack_1 : boolean;
  signal phi_stmt_2563_req_0 : boolean;
  signal phi_stmt_2813_req_1 : boolean;
  signal type_cast_2818_inst_ack_1 : boolean;
  signal type_cast_2818_inst_req_1 : boolean;
  signal phi_stmt_2556_req_1 : boolean;
  signal type_cast_2818_inst_ack_0 : boolean;
  signal type_cast_2818_inst_req_0 : boolean;
  signal type_cast_2686_inst_ack_0 : boolean;
  signal type_cast_2568_inst_req_0 : boolean;
  signal type_cast_2568_inst_ack_0 : boolean;
  signal type_cast_2568_inst_req_1 : boolean;
  signal type_cast_2568_inst_ack_1 : boolean;
  signal phi_stmt_2563_req_1 : boolean;
  signal phi_stmt_2556_ack_0 : boolean;
  signal phi_stmt_2563_ack_0 : boolean;
  signal type_cast_2686_inst_req_0 : boolean;
  signal type_cast_2617_inst_req_0 : boolean;
  signal type_cast_2617_inst_ack_0 : boolean;
  signal type_cast_2617_inst_req_1 : boolean;
  signal type_cast_2617_inst_ack_1 : boolean;
  signal phi_stmt_2614_req_0 : boolean;
  signal type_cast_2621_inst_req_0 : boolean;
  signal type_cast_2621_inst_ack_0 : boolean;
  signal type_cast_2621_inst_req_1 : boolean;
  signal type_cast_2621_inst_ack_1 : boolean;
  signal phi_stmt_2618_req_0 : boolean;
  signal phi_stmt_2614_ack_0 : boolean;
  signal phi_stmt_2618_ack_0 : boolean;
  signal type_cast_2641_inst_req_0 : boolean;
  signal type_cast_2641_inst_ack_0 : boolean;
  signal type_cast_2641_inst_req_1 : boolean;
  signal type_cast_2641_inst_ack_1 : boolean;
  signal phi_stmt_2636_req_1 : boolean;
  signal type_cast_2647_inst_req_0 : boolean;
  signal type_cast_2647_inst_ack_0 : boolean;
  signal type_cast_2647_inst_req_1 : boolean;
  signal type_cast_2647_inst_ack_1 : boolean;
  signal phi_stmt_2642_req_1 : boolean;
  signal type_cast_3391_inst_ack_0 : boolean;
  signal phi_stmt_3443_req_0 : boolean;
  signal type_cast_2639_inst_req_0 : boolean;
  signal type_cast_2639_inst_ack_0 : boolean;
  signal type_cast_2639_inst_req_1 : boolean;
  signal type_cast_2639_inst_ack_1 : boolean;
  signal phi_stmt_2636_req_0 : boolean;
  signal type_cast_2645_inst_req_0 : boolean;
  signal type_cast_2645_inst_ack_0 : boolean;
  signal type_cast_2645_inst_req_1 : boolean;
  signal type_cast_2645_inst_ack_1 : boolean;
  signal phi_stmt_2642_req_0 : boolean;
  signal phi_stmt_2636_ack_0 : boolean;
  signal phi_stmt_2642_ack_0 : boolean;
  signal phi_stmt_2683_req_1 : boolean;
  signal type_cast_2850_inst_req_0 : boolean;
  signal type_cast_2850_inst_ack_0 : boolean;
  signal type_cast_2850_inst_req_1 : boolean;
  signal type_cast_2850_inst_ack_1 : boolean;
  signal phi_stmt_2847_req_0 : boolean;
  signal type_cast_2856_inst_req_0 : boolean;
  signal type_cast_2856_inst_ack_0 : boolean;
  signal type_cast_2856_inst_req_1 : boolean;
  signal type_cast_2856_inst_ack_1 : boolean;
  signal phi_stmt_2853_req_0 : boolean;
  signal type_cast_2852_inst_req_0 : boolean;
  signal type_cast_2852_inst_ack_0 : boolean;
  signal type_cast_2852_inst_req_1 : boolean;
  signal type_cast_2852_inst_ack_1 : boolean;
  signal phi_stmt_2847_req_1 : boolean;
  signal phi_stmt_2853_req_1 : boolean;
  signal phi_stmt_2847_ack_0 : boolean;
  signal phi_stmt_2853_ack_0 : boolean;
  signal type_cast_2888_inst_req_0 : boolean;
  signal type_cast_2888_inst_ack_0 : boolean;
  signal type_cast_2888_inst_req_1 : boolean;
  signal type_cast_2888_inst_ack_1 : boolean;
  signal phi_stmt_2885_req_0 : boolean;
  signal type_cast_2892_inst_req_0 : boolean;
  signal type_cast_2892_inst_ack_0 : boolean;
  signal type_cast_2892_inst_req_1 : boolean;
  signal type_cast_2892_inst_ack_1 : boolean;
  signal phi_stmt_2889_req_0 : boolean;
  signal phi_stmt_2885_ack_0 : boolean;
  signal phi_stmt_2889_ack_0 : boolean;
  signal type_cast_2899_inst_req_0 : boolean;
  signal type_cast_2899_inst_ack_0 : boolean;
  signal type_cast_2899_inst_req_1 : boolean;
  signal type_cast_2899_inst_ack_1 : boolean;
  signal phi_stmt_2896_req_0 : boolean;
  signal phi_stmt_2902_req_0 : boolean;
  signal type_cast_2901_inst_req_0 : boolean;
  signal type_cast_2901_inst_ack_0 : boolean;
  signal type_cast_2901_inst_req_1 : boolean;
  signal type_cast_2901_inst_ack_1 : boolean;
  signal phi_stmt_2896_req_1 : boolean;
  signal type_cast_2908_inst_req_0 : boolean;
  signal type_cast_2908_inst_ack_0 : boolean;
  signal type_cast_2908_inst_req_1 : boolean;
  signal type_cast_2908_inst_ack_1 : boolean;
  signal phi_stmt_2902_req_1 : boolean;
  signal phi_stmt_2896_ack_0 : boolean;
  signal phi_stmt_2902_ack_0 : boolean;
  signal type_cast_2935_inst_req_0 : boolean;
  signal type_cast_2935_inst_ack_0 : boolean;
  signal type_cast_2935_inst_req_1 : boolean;
  signal type_cast_2935_inst_ack_1 : boolean;
  signal phi_stmt_2932_req_0 : boolean;
  signal phi_stmt_2932_ack_0 : boolean;
  signal phi_stmt_2939_req_0 : boolean;
  signal type_cast_2945_inst_req_0 : boolean;
  signal type_cast_2945_inst_ack_0 : boolean;
  signal type_cast_2945_inst_req_1 : boolean;
  signal type_cast_2945_inst_ack_1 : boolean;
  signal phi_stmt_2939_req_1 : boolean;
  signal phi_stmt_2939_ack_0 : boolean;
  signal type_cast_2954_inst_req_0 : boolean;
  signal type_cast_2954_inst_ack_0 : boolean;
  signal type_cast_2954_inst_req_1 : boolean;
  signal type_cast_2954_inst_ack_1 : boolean;
  signal phi_stmt_2949_req_1 : boolean;
  signal type_cast_2952_inst_req_0 : boolean;
  signal type_cast_2952_inst_ack_0 : boolean;
  signal type_cast_2952_inst_req_1 : boolean;
  signal type_cast_2952_inst_ack_1 : boolean;
  signal phi_stmt_2949_req_0 : boolean;
  signal phi_stmt_2949_ack_0 : boolean;
  signal type_cast_2993_inst_req_0 : boolean;
  signal type_cast_2993_inst_ack_0 : boolean;
  signal type_cast_2993_inst_req_1 : boolean;
  signal type_cast_2993_inst_ack_1 : boolean;
  signal phi_stmt_2990_req_0 : boolean;
  signal type_cast_3000_inst_req_0 : boolean;
  signal type_cast_3000_inst_ack_0 : boolean;
  signal type_cast_3000_inst_req_1 : boolean;
  signal type_cast_3000_inst_ack_1 : boolean;
  signal phi_stmt_2997_req_0 : boolean;
  signal phi_stmt_2990_req_1 : boolean;
  signal type_cast_3002_inst_req_0 : boolean;
  signal type_cast_3002_inst_ack_0 : boolean;
  signal type_cast_3002_inst_req_1 : boolean;
  signal type_cast_3002_inst_ack_1 : boolean;
  signal phi_stmt_2997_req_1 : boolean;
  signal phi_stmt_2990_ack_0 : boolean;
  signal phi_stmt_2997_ack_0 : boolean;
  signal type_cast_3051_inst_req_0 : boolean;
  signal type_cast_3051_inst_ack_0 : boolean;
  signal type_cast_3051_inst_req_1 : boolean;
  signal type_cast_3051_inst_ack_1 : boolean;
  signal phi_stmt_3048_req_0 : boolean;
  signal type_cast_3055_inst_req_0 : boolean;
  signal type_cast_3055_inst_ack_0 : boolean;
  signal type_cast_3055_inst_req_1 : boolean;
  signal type_cast_3055_inst_ack_1 : boolean;
  signal phi_stmt_3052_req_0 : boolean;
  signal phi_stmt_3048_ack_0 : boolean;
  signal phi_stmt_3052_ack_0 : boolean;
  signal type_cast_3080_inst_req_0 : boolean;
  signal type_cast_3080_inst_ack_0 : boolean;
  signal type_cast_3080_inst_req_1 : boolean;
  signal type_cast_3080_inst_ack_1 : boolean;
  signal phi_stmt_3075_req_1 : boolean;
  signal type_cast_3086_inst_req_0 : boolean;
  signal type_cast_3086_inst_ack_0 : boolean;
  signal type_cast_3086_inst_req_1 : boolean;
  signal type_cast_3086_inst_ack_1 : boolean;
  signal phi_stmt_3081_req_1 : boolean;
  signal type_cast_3078_inst_req_0 : boolean;
  signal type_cast_3078_inst_ack_0 : boolean;
  signal type_cast_3078_inst_req_1 : boolean;
  signal type_cast_3078_inst_ack_1 : boolean;
  signal phi_stmt_3075_req_0 : boolean;
  signal type_cast_3084_inst_req_0 : boolean;
  signal type_cast_3084_inst_ack_0 : boolean;
  signal type_cast_3084_inst_req_1 : boolean;
  signal type_cast_3084_inst_ack_1 : boolean;
  signal phi_stmt_3081_req_0 : boolean;
  signal phi_stmt_3075_ack_0 : boolean;
  signal phi_stmt_3081_ack_0 : boolean;
  signal phi_stmt_3122_req_1 : boolean;
  signal type_cast_3125_inst_req_0 : boolean;
  signal type_cast_3125_inst_ack_0 : boolean;
  signal type_cast_3125_inst_req_1 : boolean;
  signal type_cast_3125_inst_ack_1 : boolean;
  signal phi_stmt_3122_req_0 : boolean;
  signal phi_stmt_3122_ack_0 : boolean;
  signal type_cast_3391_inst_req_0 : boolean;
  signal type_cast_3446_inst_ack_1 : boolean;
  signal type_cast_3446_inst_req_1 : boolean;
  signal type_cast_3264_inst_req_0 : boolean;
  signal type_cast_3264_inst_ack_0 : boolean;
  signal type_cast_3264_inst_req_1 : boolean;
  signal type_cast_3264_inst_ack_1 : boolean;
  signal phi_stmt_3259_req_1 : boolean;
  signal type_cast_3446_inst_ack_0 : boolean;
  signal type_cast_3446_inst_req_0 : boolean;
  signal phi_stmt_3265_req_1 : boolean;
  signal type_cast_3262_inst_req_0 : boolean;
  signal type_cast_3262_inst_ack_0 : boolean;
  signal type_cast_3262_inst_req_1 : boolean;
  signal type_cast_3262_inst_ack_1 : boolean;
  signal phi_stmt_3259_req_0 : boolean;
  signal type_cast_3268_inst_req_0 : boolean;
  signal type_cast_3268_inst_ack_0 : boolean;
  signal type_cast_3268_inst_req_1 : boolean;
  signal type_cast_3268_inst_ack_1 : boolean;
  signal phi_stmt_3265_req_0 : boolean;
  signal phi_stmt_3259_ack_0 : boolean;
  signal phi_stmt_3265_ack_0 : boolean;
  signal type_cast_3391_inst_req_1 : boolean;
  signal phi_stmt_3395_ack_0 : boolean;
  signal type_cast_3296_inst_req_0 : boolean;
  signal type_cast_3296_inst_ack_0 : boolean;
  signal type_cast_3296_inst_req_1 : boolean;
  signal type_cast_3296_inst_ack_1 : boolean;
  signal phi_stmt_3395_req_0 : boolean;
  signal phi_stmt_3293_req_0 : boolean;
  signal type_cast_3302_inst_req_0 : boolean;
  signal type_cast_3302_inst_ack_0 : boolean;
  signal type_cast_3302_inst_req_1 : boolean;
  signal type_cast_3302_inst_ack_1 : boolean;
  signal phi_stmt_3299_req_0 : boolean;
  signal type_cast_3398_inst_ack_1 : boolean;
  signal type_cast_3398_inst_req_1 : boolean;
  signal type_cast_3298_inst_req_0 : boolean;
  signal type_cast_3298_inst_ack_0 : boolean;
  signal type_cast_3298_inst_req_1 : boolean;
  signal type_cast_3298_inst_ack_1 : boolean;
  signal phi_stmt_3293_req_1 : boolean;
  signal type_cast_3398_inst_ack_0 : boolean;
  signal type_cast_3398_inst_req_0 : boolean;
  signal phi_stmt_3299_req_1 : boolean;
  signal phi_stmt_3293_ack_0 : boolean;
  signal phi_stmt_3299_ack_0 : boolean;
  signal phi_stmt_3385_req_0 : boolean;
  signal type_cast_3338_inst_req_0 : boolean;
  signal type_cast_3338_inst_ack_0 : boolean;
  signal type_cast_3338_inst_req_1 : boolean;
  signal type_cast_3338_inst_ack_1 : boolean;
  signal phi_stmt_3335_req_0 : boolean;
  signal phi_stmt_3395_req_1 : boolean;
  signal type_cast_3334_inst_req_0 : boolean;
  signal type_cast_3334_inst_ack_0 : boolean;
  signal type_cast_3400_inst_ack_1 : boolean;
  signal type_cast_3334_inst_req_1 : boolean;
  signal type_cast_3334_inst_ack_1 : boolean;
  signal phi_stmt_3331_req_0 : boolean;
  signal phi_stmt_3331_ack_0 : boolean;
  signal phi_stmt_3335_ack_0 : boolean;
  signal type_cast_3400_inst_req_1 : boolean;
  signal type_cast_3400_inst_ack_0 : boolean;
  signal type_cast_3400_inst_req_0 : boolean;
  signal phi_stmt_3348_req_0 : boolean;
  signal type_cast_3345_inst_req_0 : boolean;
  signal type_cast_3345_inst_ack_0 : boolean;
  signal type_cast_3345_inst_req_1 : boolean;
  signal type_cast_3345_inst_ack_1 : boolean;
  signal phi_stmt_3342_req_0 : boolean;
  signal type_cast_3354_inst_req_0 : boolean;
  signal type_cast_3354_inst_ack_0 : boolean;
  signal type_cast_3354_inst_req_1 : boolean;
  signal type_cast_3354_inst_ack_1 : boolean;
  signal phi_stmt_3348_req_1 : boolean;
  signal type_cast_3347_inst_req_0 : boolean;
  signal type_cast_3347_inst_ack_0 : boolean;
  signal type_cast_3347_inst_req_1 : boolean;
  signal type_cast_3347_inst_ack_1 : boolean;
  signal phi_stmt_3342_req_1 : boolean;
  signal phi_stmt_3342_ack_0 : boolean;
  signal phi_stmt_3348_ack_0 : boolean;
  signal phi_stmt_3385_ack_0 : boolean;
  signal phi_stmt_3385_req_1 : boolean;
  signal type_cast_3381_inst_req_0 : boolean;
  signal type_cast_3381_inst_ack_0 : boolean;
  signal type_cast_3391_inst_ack_1 : boolean;
  signal type_cast_3381_inst_req_1 : boolean;
  signal type_cast_3381_inst_ack_1 : boolean;
  signal phi_stmt_3378_req_0 : boolean;
  signal phi_stmt_3378_ack_0 : boolean;
  signal type_cast_3439_inst_req_0 : boolean;
  signal type_cast_3439_inst_ack_0 : boolean;
  signal type_cast_3439_inst_req_1 : boolean;
  signal type_cast_3439_inst_ack_1 : boolean;
  signal phi_stmt_3436_req_0 : boolean;
  signal type_cast_3448_inst_req_0 : boolean;
  signal type_cast_3448_inst_ack_0 : boolean;
  signal type_cast_3448_inst_req_1 : boolean;
  signal type_cast_3448_inst_ack_1 : boolean;
  signal phi_stmt_3443_req_1 : boolean;
  signal phi_stmt_3436_req_1 : boolean;
  signal phi_stmt_3436_ack_0 : boolean;
  signal phi_stmt_3443_ack_0 : boolean;
  signal type_cast_3501_inst_req_0 : boolean;
  signal type_cast_3501_inst_ack_0 : boolean;
  signal type_cast_3501_inst_req_1 : boolean;
  signal type_cast_3501_inst_ack_1 : boolean;
  signal phi_stmt_3498_req_0 : boolean;
  signal type_cast_3497_inst_req_0 : boolean;
  signal type_cast_3497_inst_ack_0 : boolean;
  signal type_cast_3497_inst_req_1 : boolean;
  signal type_cast_3497_inst_ack_1 : boolean;
  signal phi_stmt_3494_req_0 : boolean;
  signal phi_stmt_3494_ack_0 : boolean;
  signal phi_stmt_3498_ack_0 : boolean;
  signal type_cast_3526_inst_req_0 : boolean;
  signal type_cast_3526_inst_ack_0 : boolean;
  signal type_cast_3526_inst_req_1 : boolean;
  signal type_cast_3526_inst_ack_1 : boolean;
  signal phi_stmt_3521_req_1 : boolean;
  signal type_cast_3532_inst_req_0 : boolean;
  signal type_cast_3532_inst_ack_0 : boolean;
  signal type_cast_3532_inst_req_1 : boolean;
  signal type_cast_3532_inst_ack_1 : boolean;
  signal phi_stmt_3527_req_1 : boolean;
  signal type_cast_3524_inst_req_0 : boolean;
  signal type_cast_3524_inst_ack_0 : boolean;
  signal type_cast_3524_inst_req_1 : boolean;
  signal type_cast_3524_inst_ack_1 : boolean;
  signal phi_stmt_3521_req_0 : boolean;
  signal type_cast_3530_inst_req_0 : boolean;
  signal type_cast_3530_inst_ack_0 : boolean;
  signal type_cast_3530_inst_req_1 : boolean;
  signal type_cast_3530_inst_ack_1 : boolean;
  signal phi_stmt_3527_req_0 : boolean;
  signal phi_stmt_3521_ack_0 : boolean;
  signal phi_stmt_3527_ack_0 : boolean;
  signal phi_stmt_3568_req_1 : boolean;
  signal type_cast_3571_inst_req_0 : boolean;
  signal type_cast_3571_inst_ack_0 : boolean;
  signal type_cast_3571_inst_req_1 : boolean;
  signal type_cast_3571_inst_ack_1 : boolean;
  signal phi_stmt_3568_req_0 : boolean;
  signal phi_stmt_3568_ack_0 : boolean;
  signal phi_stmt_3626_req_2 : boolean;
  signal type_cast_3629_inst_req_0 : boolean;
  signal type_cast_3629_inst_ack_0 : boolean;
  signal type_cast_3629_inst_req_1 : boolean;
  signal type_cast_3629_inst_ack_1 : boolean;
  signal phi_stmt_3626_req_0 : boolean;
  signal phi_stmt_3626_req_1 : boolean;
  signal phi_stmt_3626_ack_0 : boolean;
  signal phi_stmt_3687_req_1 : boolean;
  signal phi_stmt_3687_req_2 : boolean;
  signal type_cast_3690_inst_req_0 : boolean;
  signal type_cast_3690_inst_ack_0 : boolean;
  signal type_cast_3690_inst_req_1 : boolean;
  signal type_cast_3690_inst_ack_1 : boolean;
  signal phi_stmt_3687_req_0 : boolean;
  signal phi_stmt_3687_ack_0 : boolean;
  signal type_cast_3725_inst_req_0 : boolean;
  signal type_cast_3725_inst_ack_0 : boolean;
  signal type_cast_3725_inst_req_1 : boolean;
  signal type_cast_3725_inst_ack_1 : boolean;
  signal phi_stmt_3722_req_0 : boolean;
  signal type_cast_3731_inst_req_0 : boolean;
  signal type_cast_3731_inst_ack_0 : boolean;
  signal type_cast_3731_inst_req_1 : boolean;
  signal type_cast_3731_inst_ack_1 : boolean;
  signal phi_stmt_3728_req_0 : boolean;
  signal type_cast_3727_inst_req_0 : boolean;
  signal type_cast_3727_inst_ack_0 : boolean;
  signal type_cast_3727_inst_req_1 : boolean;
  signal type_cast_3727_inst_ack_1 : boolean;
  signal phi_stmt_3722_req_1 : boolean;
  signal phi_stmt_3728_req_1 : boolean;
  signal phi_stmt_3722_ack_0 : boolean;
  signal phi_stmt_3728_ack_0 : boolean;
  signal type_cast_3760_inst_req_0 : boolean;
  signal type_cast_3760_inst_ack_0 : boolean;
  signal type_cast_3760_inst_req_1 : boolean;
  signal type_cast_3760_inst_ack_1 : boolean;
  signal phi_stmt_3757_req_0 : boolean;
  signal type_cast_3767_inst_req_0 : boolean;
  signal type_cast_3767_inst_ack_0 : boolean;
  signal type_cast_3767_inst_req_1 : boolean;
  signal type_cast_3767_inst_ack_1 : boolean;
  signal phi_stmt_3764_req_0 : boolean;
  signal phi_stmt_3757_req_1 : boolean;
  signal phi_stmt_3764_req_1 : boolean;
  signal phi_stmt_3757_ack_0 : boolean;
  signal phi_stmt_3764_ack_0 : boolean;
  signal type_cast_3799_inst_req_0 : boolean;
  signal type_cast_3799_inst_ack_0 : boolean;
  signal type_cast_3799_inst_req_1 : boolean;
  signal type_cast_3799_inst_ack_1 : boolean;
  signal phi_stmt_3796_req_0 : boolean;
  signal type_cast_3803_inst_req_0 : boolean;
  signal type_cast_3803_inst_ack_0 : boolean;
  signal type_cast_3803_inst_req_1 : boolean;
  signal type_cast_3803_inst_ack_1 : boolean;
  signal phi_stmt_3800_req_0 : boolean;
  signal phi_stmt_3796_ack_0 : boolean;
  signal phi_stmt_3800_ack_0 : boolean;
  signal phi_stmt_3807_req_0 : boolean;
  signal phi_stmt_3814_req_0 : boolean;
  signal type_cast_3813_inst_req_0 : boolean;
  signal type_cast_3813_inst_ack_0 : boolean;
  signal type_cast_3813_inst_req_1 : boolean;
  signal type_cast_3813_inst_ack_1 : boolean;
  signal phi_stmt_3807_req_1 : boolean;
  signal type_cast_3820_inst_req_0 : boolean;
  signal type_cast_3820_inst_ack_0 : boolean;
  signal type_cast_3820_inst_req_1 : boolean;
  signal type_cast_3820_inst_ack_1 : boolean;
  signal phi_stmt_3814_req_1 : boolean;
  signal phi_stmt_3807_ack_0 : boolean;
  signal phi_stmt_3814_ack_0 : boolean;
  signal type_cast_3848_inst_req_0 : boolean;
  signal type_cast_3848_inst_ack_0 : boolean;
  signal type_cast_3848_inst_req_1 : boolean;
  signal type_cast_3848_inst_ack_1 : boolean;
  signal phi_stmt_3845_req_0 : boolean;
  signal phi_stmt_3845_ack_0 : boolean;
  signal type_cast_3911_inst_req_0 : boolean;
  signal type_cast_3911_inst_ack_0 : boolean;
  signal type_cast_3911_inst_req_1 : boolean;
  signal type_cast_3911_inst_ack_1 : boolean;
  signal phi_stmt_3908_req_0 : boolean;
  signal type_cast_3918_inst_req_0 : boolean;
  signal type_cast_3918_inst_ack_0 : boolean;
  signal type_cast_3918_inst_req_1 : boolean;
  signal type_cast_3918_inst_ack_1 : boolean;
  signal phi_stmt_3915_req_0 : boolean;
  signal phi_stmt_3908_req_1 : boolean;
  signal type_cast_3920_inst_req_0 : boolean;
  signal type_cast_3920_inst_ack_0 : boolean;
  signal type_cast_3920_inst_req_1 : boolean;
  signal type_cast_3920_inst_ack_1 : boolean;
  signal phi_stmt_3915_req_1 : boolean;
  signal phi_stmt_3908_ack_0 : boolean;
  signal phi_stmt_3915_ack_0 : boolean;
  signal type_cast_3969_inst_req_0 : boolean;
  signal type_cast_3969_inst_ack_0 : boolean;
  signal type_cast_3969_inst_req_1 : boolean;
  signal type_cast_3969_inst_ack_1 : boolean;
  signal phi_stmt_3966_req_0 : boolean;
  signal type_cast_3973_inst_req_0 : boolean;
  signal type_cast_3973_inst_ack_0 : boolean;
  signal type_cast_3973_inst_req_1 : boolean;
  signal type_cast_3973_inst_ack_1 : boolean;
  signal phi_stmt_3970_req_0 : boolean;
  signal phi_stmt_3966_ack_0 : boolean;
  signal phi_stmt_3970_ack_0 : boolean;
  signal type_cast_3993_inst_req_0 : boolean;
  signal type_cast_3993_inst_ack_0 : boolean;
  signal type_cast_3993_inst_req_1 : boolean;
  signal type_cast_3993_inst_ack_1 : boolean;
  signal phi_stmt_3988_req_1 : boolean;
  signal type_cast_3999_inst_req_0 : boolean;
  signal type_cast_3999_inst_ack_0 : boolean;
  signal type_cast_3999_inst_req_1 : boolean;
  signal type_cast_3999_inst_ack_1 : boolean;
  signal phi_stmt_3994_req_1 : boolean;
  signal type_cast_3991_inst_req_0 : boolean;
  signal type_cast_3991_inst_ack_0 : boolean;
  signal type_cast_3991_inst_req_1 : boolean;
  signal type_cast_3991_inst_ack_1 : boolean;
  signal phi_stmt_3988_req_0 : boolean;
  signal type_cast_3997_inst_req_0 : boolean;
  signal type_cast_3997_inst_ack_0 : boolean;
  signal type_cast_3997_inst_req_1 : boolean;
  signal type_cast_3997_inst_ack_1 : boolean;
  signal phi_stmt_3994_req_0 : boolean;
  signal phi_stmt_3988_ack_0 : boolean;
  signal phi_stmt_3994_ack_0 : boolean;
  signal phi_stmt_4035_req_1 : boolean;
  signal type_cast_4038_inst_req_0 : boolean;
  signal type_cast_4038_inst_ack_0 : boolean;
  signal type_cast_4038_inst_req_1 : boolean;
  signal type_cast_4038_inst_ack_1 : boolean;
  signal phi_stmt_4035_req_0 : boolean;
  signal phi_stmt_4035_ack_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "vector_control_daemon_input_buffer", -- 
      buffer_size => 1,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  vector_control_daemon_CP_10259_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "vector_control_daemon_out_buffer", -- 
      buffer_size => 1,
      data_width => tag_length + 0, 
      kill_counter_range => 1) -- 
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      kill => default_zero_sig,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= vector_control_daemon_CP_10259_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= vector_control_daemon_CP_10259_start & tag_ilock_write_ack_symbol;
    gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= vector_control_daemon_CP_10259_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  vector_control_daemon_CP_10259: Block -- control-path 
    signal cp_elements: BooleanArray(2585 downto 0);
    -- 
  begin -- 
    cp_elements(0) <= vector_control_daemon_CP_10259_start;
    vector_control_daemon_CP_10259_symbol <= cp_elements(1);
    -- CP-element group 0 transition  place  bypass 
    -- predecessors 
    -- successors 1277 
    -- members (4) 
      -- 	$entry
      -- 	branch_block_stmt_2042/$entry
      -- 	branch_block_stmt_2042/branch_block_stmt_2042__entry__
      -- 	branch_block_stmt_2042/bb_0_bb_1
      -- 
    -- CP-element group 1 transition  place  bypass 
    -- predecessors 
    -- successors 
    -- members (3) 
      -- 	$exit
      -- 	branch_block_stmt_2042/$exit
      -- 	branch_block_stmt_2042/branch_block_stmt_2042__exit__
      -- 
    cp_elements(1) <= false; 
    -- CP-element group 2 place  bypass 
    -- predecessors 1316 
    -- successors 79 
    -- members (2) 
      -- 	branch_block_stmt_2042/merge_stmt_2044__exit__
      -- 	branch_block_stmt_2042/assign_stmt_2069__entry__
      -- 
    cp_elements(2) <= cp_elements(1316);
    -- CP-element group 3 merge  place  bypass 
    -- predecessors 123 129 
    -- successors 130 
    -- members (2) 
      -- 	branch_block_stmt_2042/merge_stmt_2118__exit__
      -- 	branch_block_stmt_2042/assign_stmt_2124__entry__
      -- 
    cp_elements(3) <= OrReduce(cp_elements(123) & cp_elements(129));
    -- CP-element group 4 merge  fork  transition  place  bypass 
    -- predecessors 135 141 
    -- successors 1323 1325 
    -- members (7) 
      -- 	branch_block_stmt_2042/merge_stmt_2131__exit__
      -- 	branch_block_stmt_2042/bb_3_bb_4
      -- 	branch_block_stmt_2042/bb_3_bb_4_PhiReq/$entry
      -- 	branch_block_stmt_2042/bb_3_bb_4_PhiReq/phi_stmt_2134/$entry
      -- 	branch_block_stmt_2042/bb_3_bb_4_PhiReq/phi_stmt_2134/phi_stmt_2134_sources/$entry
      -- 	branch_block_stmt_2042/bb_3_bb_4_PhiReq/phi_stmt_2134/phi_stmt_2134_sources/type_cast_2137/$entry
      -- 	branch_block_stmt_2042/bb_3_bb_4_PhiReq/phi_stmt_2134/phi_stmt_2134_sources/type_cast_2137/SplitProtocol/$entry
      -- 
    cp_elements(4) <= OrReduce(cp_elements(135) & cp_elements(141));
    -- CP-element group 5 merge  place  bypass 
    -- predecessors 155 161 
    -- successors 162 
    -- members (2) 
      -- 	branch_block_stmt_2042/merge_stmt_2168__exit__
      -- 	branch_block_stmt_2042/assign_stmt_2174__entry__
      -- 
    cp_elements(5) <= OrReduce(cp_elements(155) & cp_elements(161));
    -- CP-element group 6 merge  place  bypass 
    -- predecessors 167 173 
    -- successors 174 
    -- members (2) 
      -- 	branch_block_stmt_2042/merge_stmt_2181__exit__
      -- 	branch_block_stmt_2042/assign_stmt_2187__entry__
      -- 
    cp_elements(6) <= OrReduce(cp_elements(167) & cp_elements(173));
    -- CP-element group 7 merge  place  bypass 
    -- predecessors 187 191 
    -- successors 194 
    -- members (2) 
      -- 	branch_block_stmt_2042/merge_stmt_2217__exit__
      -- 	branch_block_stmt_2042/assign_stmt_2223__entry__
      -- 
    cp_elements(7) <= OrReduce(cp_elements(187) & cp_elements(191));
    -- CP-element group 8 merge  place  bypass 
    -- predecessors 199 205 
    -- successors 206 
    -- members (2) 
      -- 	branch_block_stmt_2042/merge_stmt_2230__exit__
      -- 	branch_block_stmt_2042/assign_stmt_2236_to_assign_stmt_2248__entry__
      -- 
    cp_elements(8) <= OrReduce(cp_elements(199) & cp_elements(205));
    -- CP-element group 9 merge  place  bypass 
    -- predecessors 222 228 
    -- successors 229 
    -- members (2) 
      -- 	branch_block_stmt_2042/merge_stmt_2263__exit__
      -- 	branch_block_stmt_2042/assign_stmt_2269_to_assign_stmt_2281__entry__
      -- 
    cp_elements(9) <= OrReduce(cp_elements(222) & cp_elements(228));
    -- CP-element group 10 branch  place  bypass 
    -- predecessors 272 
    -- successors 273 274 
    -- members (2) 
      -- 	branch_block_stmt_2042/assign_stmt_2321_to_assign_stmt_2342__exit__
      -- 	branch_block_stmt_2042/if_stmt_2343__entry__
      -- 
    cp_elements(10) <= cp_elements(272);
    -- CP-element group 11 merge  place  bypass 
    -- predecessors 273 279 
    -- successors 280 
    -- members (2) 
      -- 	branch_block_stmt_2042/merge_stmt_2349__exit__
      -- 	branch_block_stmt_2042/assign_stmt_2355_to_assign_stmt_2367__entry__
      -- 
    cp_elements(11) <= OrReduce(cp_elements(273) & cp_elements(279));
    -- CP-element group 12 place  bypass 
    -- predecessors 1448 
    -- successors 291 
    -- members (2) 
      -- 	branch_block_stmt_2042/merge_stmt_2369__exit__
      -- 	branch_block_stmt_2042/assign_stmt_2389_to_assign_stmt_2395__entry__
      -- 
    cp_elements(12) <= cp_elements(1448);
    -- CP-element group 13 merge  place  bypass 
    -- predecessors 299 303 
    -- successors 1463 
    -- members (2) 
      -- 	branch_block_stmt_2042/merge_stmt_2402__exit__
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi36x_xpreheader_bbx_xnphx_xix_xix_xi36
      -- 
    cp_elements(13) <= OrReduce(cp_elements(299) & cp_elements(303));
    -- CP-element group 14 place  bypass 
    -- predecessors 1477 
    -- successors 306 
    -- members (2) 
      -- 	branch_block_stmt_2042/merge_stmt_2404__exit__
      -- 	branch_block_stmt_2042/assign_stmt_2425_to_assign_stmt_2436__entry__
      -- 
    cp_elements(14) <= cp_elements(1477);
    -- CP-element group 15 branch  place  bypass 
    -- predecessors 320 
    -- successors 321 322 
    -- members (2) 
      -- 	branch_block_stmt_2042/assign_stmt_2425_to_assign_stmt_2436__exit__
      -- 	branch_block_stmt_2042/if_stmt_2437__entry__
      -- 
    cp_elements(15) <= cp_elements(320);
    -- CP-element group 16 merge  place  bypass 
    -- predecessors 321 1496 
    -- successors 1507 
    -- members (2) 
      -- 	branch_block_stmt_2042/merge_stmt_2443__exit__
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi39x_xloopexit_xx_x_crit_edgex_xix_xix_xi39
      -- 
    cp_elements(16) <= OrReduce(cp_elements(321) & cp_elements(1496));
    -- CP-element group 17 place  bypass 
    -- predecessors 1525 
    -- successors 328 
    -- members (2) 
      -- 	branch_block_stmt_2042/merge_stmt_2454__exit__
      -- 	branch_block_stmt_2042/assign_stmt_2474_to_assign_stmt_2485__entry__
      -- 
    cp_elements(17) <= cp_elements(1525);
    -- CP-element group 18 branch  place  bypass 
    -- predecessors 344 
    -- successors 345 346 
    -- members (2) 
      -- 	branch_block_stmt_2042/assign_stmt_2474_to_assign_stmt_2485__exit__
      -- 	branch_block_stmt_2042/if_stmt_2486__entry__
      -- 
    cp_elements(18) <= cp_elements(344);
    -- CP-element group 19 merge  place  bypass 
    -- predecessors 345 1531 
    -- successors 352 
    -- members (2) 
      -- 	branch_block_stmt_2042/merge_stmt_2492__exit__
      -- 	branch_block_stmt_2042/assign_stmt_2503_to_assign_stmt_2546__entry__
      -- 
    cp_elements(19) <= OrReduce(cp_elements(345) & cp_elements(1531));
    -- CP-element group 20 branch  place  bypass 
    -- predecessors 384 
    -- successors 385 386 
    -- members (2) 
      -- 	branch_block_stmt_2042/assign_stmt_2503_to_assign_stmt_2546__exit__
      -- 	branch_block_stmt_2042/if_stmt_2547__entry__
      -- 
    cp_elements(20) <= cp_elements(384);
    -- CP-element group 21 merge  place  bypass 
    -- predecessors 385 389 
    -- successors 1552 
    -- members (2) 
      -- 	branch_block_stmt_2042/merge_stmt_2553__exit__
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi45x_xpreheader_udiv32x_xexitx_xix_xi45
      -- 
    cp_elements(21) <= OrReduce(cp_elements(385) & cp_elements(389));
    -- CP-element group 22 place  bypass 
    -- predecessors 1574 
    -- successors 392 
    -- members (2) 
      -- 	branch_block_stmt_2042/merge_stmt_2555__exit__
      -- 	branch_block_stmt_2042/assign_stmt_2575_to_assign_stmt_2606__entry__
      -- 
    cp_elements(22) <= cp_elements(1574);
    -- CP-element group 23 branch  place  bypass 
    -- predecessors 418 
    -- successors 419 420 
    -- members (2) 
      -- 	branch_block_stmt_2042/assign_stmt_2575_to_assign_stmt_2606__exit__
      -- 	branch_block_stmt_2042/if_stmt_2607__entry__
      -- 
    cp_elements(23) <= cp_elements(418);
    -- CP-element group 24 merge  place  bypass 
    -- predecessors 419 1593 
    -- successors 426 
    -- members (2) 
      -- 	branch_block_stmt_2042/merge_stmt_2613__exit__
      -- 	branch_block_stmt_2042/assign_stmt_2628_to_assign_stmt_2633__entry__
      -- 
    cp_elements(24) <= OrReduce(cp_elements(419) & cp_elements(1593));
    -- CP-element group 25 place  bypass 
    -- predecessors 1650 
    -- successors 436 
    -- members (2) 
      -- 	branch_block_stmt_2042/merge_stmt_2635__exit__
      -- 	branch_block_stmt_2042/assign_stmt_2654_to_assign_stmt_2680__entry__
      -- 
    cp_elements(25) <= cp_elements(1650);
    -- CP-element group 26 branch  place  bypass 
    -- predecessors 480 
    -- successors 481 482 
    -- members (2) 
      -- 	branch_block_stmt_2042/assign_stmt_2696_to_assign_stmt_2716__exit__
      -- 	branch_block_stmt_2042/if_stmt_2717__entry__
      -- 
    cp_elements(26) <= cp_elements(480);
    -- CP-element group 27 merge  place  bypass 
    -- predecessors 481 487 
    -- successors 488 
    -- members (2) 
      -- 	branch_block_stmt_2042/assign_stmt_2729_to_assign_stmt_2799__entry__
      -- 	branch_block_stmt_2042/merge_stmt_2723__exit__
      -- 
    cp_elements(27) <= OrReduce(cp_elements(481) & cp_elements(487));
    -- CP-element group 28 branch  place  bypass 
    -- predecessors 536 
    -- successors 537 538 
    -- members (2) 
      -- 	branch_block_stmt_2042/assign_stmt_2729_to_assign_stmt_2799__exit__
      -- 	branch_block_stmt_2042/switch_stmt_2800__entry__
      -- 
    cp_elements(28) <= cp_elements(536);
    -- CP-element group 29 merge  place  bypass 
    -- predecessors 537 559 
    -- successors 1662 
    -- members (2) 
      -- 	branch_block_stmt_2042/merge_stmt_2810__exit__
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xix_xi5x_xpreheader_bbx_xnph7x_xix_xix_xi5
      -- 
    cp_elements(29) <= OrReduce(cp_elements(537) & cp_elements(559));
    -- CP-element group 30 place  bypass 
    -- predecessors 1704 
    -- successors 560 
    -- members (2) 
      -- 	branch_block_stmt_2042/merge_stmt_2812__exit__
      -- 	branch_block_stmt_2042/assign_stmt_2832_to_assign_stmt_2837__entry__
      -- 
    cp_elements(30) <= cp_elements(1704);
    -- CP-element group 31 merge  place  bypass 
    -- predecessors 570 574 
    -- successors 1725 
    -- members (2) 
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi8x_xpreheader_bbx_xnphx_xix_xix_xi8
      -- 	branch_block_stmt_2042/merge_stmt_2844__exit__
      -- 
    cp_elements(31) <= OrReduce(cp_elements(570) & cp_elements(574));
    -- CP-element group 32 place  bypass 
    -- predecessors 1747 
    -- successors 577 
    -- members (2) 
      -- 	branch_block_stmt_2042/merge_stmt_2846__exit__
      -- 	branch_block_stmt_2042/assign_stmt_2866_to_assign_stmt_2877__entry__
      -- 
    cp_elements(32) <= cp_elements(1747);
    -- CP-element group 33 branch  place  bypass 
    -- predecessors 591 
    -- successors 592 593 
    -- members (2) 
      -- 	branch_block_stmt_2042/assign_stmt_2866_to_assign_stmt_2877__exit__
      -- 	branch_block_stmt_2042/if_stmt_2878__entry__
      -- 
    cp_elements(33) <= cp_elements(591);
    -- CP-element group 34 merge  place  bypass 
    -- predecessors 592 1766 
    -- successors 1785 
    -- members (2) 
      -- 	branch_block_stmt_2042/merge_stmt_2884__exit__
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi11x_xloopexit_xx_x_crit_edgex_xix_xix_xi11
      -- 
    cp_elements(34) <= OrReduce(cp_elements(592) & cp_elements(1766));
    -- CP-element group 35 place  bypass 
    -- predecessors 1809 
    -- successors 599 
    -- members (2) 
      -- 	branch_block_stmt_2042/merge_stmt_2895__exit__
      -- 	branch_block_stmt_2042/assign_stmt_2914_to_assign_stmt_2924__entry__
      -- 
    cp_elements(35) <= cp_elements(1809);
    -- CP-element group 36 branch  place  bypass 
    -- predecessors 617 
    -- successors 618 619 
    -- members (2) 
      -- 	branch_block_stmt_2042/if_stmt_2925__entry__
      -- 	branch_block_stmt_2042/assign_stmt_2914_to_assign_stmt_2924__exit__
      -- 
    cp_elements(36) <= cp_elements(617);
    -- CP-element group 37 merge  fork  transition  place  bypass 
    -- predecessors 618 1815 
    -- successors 1819 1821 
    -- members (7) 
      -- 	branch_block_stmt_2042/xx_xloopexitx_xix_xix_xi13x_xloopexit_xx_xloopexitx_xix_xix_xi13
      -- 	branch_block_stmt_2042/merge_stmt_2931__exit__
      -- 	branch_block_stmt_2042/xx_xloopexitx_xix_xix_xi13x_xloopexit_xx_xloopexitx_xix_xix_xi13_PhiReq/$entry
      -- 	branch_block_stmt_2042/xx_xloopexitx_xix_xix_xi13x_xloopexit_xx_xloopexitx_xix_xix_xi13_PhiReq/phi_stmt_2939/$entry
      -- 	branch_block_stmt_2042/xx_xloopexitx_xix_xix_xi13x_xloopexit_xx_xloopexitx_xix_xix_xi13_PhiReq/phi_stmt_2939/phi_stmt_2939_sources/$entry
      -- 	branch_block_stmt_2042/xx_xloopexitx_xix_xix_xi13x_xloopexit_xx_xloopexitx_xix_xix_xi13_PhiReq/phi_stmt_2939/phi_stmt_2939_sources/type_cast_2945/$entry
      -- 	branch_block_stmt_2042/xx_xloopexitx_xix_xix_xi13x_xloopexit_xx_xloopexitx_xix_xix_xi13_PhiReq/phi_stmt_2939/phi_stmt_2939_sources/type_cast_2945/SplitProtocol/$entry
      -- 
    cp_elements(37) <= OrReduce(cp_elements(618) & cp_elements(1815));
    -- CP-element group 38 merge  place  bypass 
    -- predecessors 643 647 
    -- successors 1872 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi20x_xpreheader_udiv32x_xexitx_xix_xi20
      -- 	branch_block_stmt_2042/merge_stmt_2987__exit__
      -- 
    cp_elements(38) <= OrReduce(cp_elements(643) & cp_elements(647));
    -- CP-element group 39 place  bypass 
    -- predecessors 1894 
    -- successors 650 
    -- members (2) 
      -- 	branch_block_stmt_2042/assign_stmt_3009_to_assign_stmt_3040__entry__
      -- 	branch_block_stmt_2042/merge_stmt_2989__exit__
      -- 
    cp_elements(39) <= cp_elements(1894);
    -- CP-element group 40 branch  place  bypass 
    -- predecessors 676 
    -- successors 677 678 
    -- members (2) 
      -- 	branch_block_stmt_2042/if_stmt_3041__entry__
      -- 	branch_block_stmt_2042/assign_stmt_3009_to_assign_stmt_3040__exit__
      -- 
    cp_elements(40) <= cp_elements(676);
    -- CP-element group 41 merge  place  bypass 
    -- predecessors 677 1913 
    -- successors 684 
    -- members (2) 
      -- 	branch_block_stmt_2042/assign_stmt_3062_to_assign_stmt_3072__entry__
      -- 	branch_block_stmt_2042/merge_stmt_3047__exit__
      -- 
    cp_elements(41) <= OrReduce(cp_elements(677) & cp_elements(1913));
    -- CP-element group 42 place  bypass 
    -- predecessors 1970 
    -- successors 699 
    -- members (2) 
      -- 	branch_block_stmt_2042/assign_stmt_3093_to_assign_stmt_3119__entry__
      -- 	branch_block_stmt_2042/merge_stmt_3074__exit__
      -- 
    cp_elements(42) <= cp_elements(1970);
    -- CP-element group 43 branch  place  bypass 
    -- predecessors 747 
    -- successors 748 749 
    -- members (2) 
      -- 	branch_block_stmt_2042/if_stmt_3163__entry__
      -- 	branch_block_stmt_2042/assign_stmt_3135_to_assign_stmt_3162__exit__
      -- 
    cp_elements(43) <= cp_elements(747);
    -- CP-element group 44 merge  place  bypass 
    -- predecessors 748 754 
    -- successors 755 
    -- members (2) 
      -- 	branch_block_stmt_2042/assign_stmt_3175_to_assign_stmt_3245__entry__
      -- 	branch_block_stmt_2042/merge_stmt_3169__exit__
      -- 
    cp_elements(44) <= OrReduce(cp_elements(748) & cp_elements(754));
    -- CP-element group 45 branch  place  bypass 
    -- predecessors 803 
    -- successors 804 805 
    -- members (2) 
      -- 	branch_block_stmt_2042/switch_stmt_3246__entry__
      -- 	branch_block_stmt_2042/assign_stmt_3175_to_assign_stmt_3245__exit__
      -- 
    cp_elements(45) <= cp_elements(803);
    -- CP-element group 46 merge  place  bypass 
    -- predecessors 804 826 
    -- successors 1982 
    -- members (2) 
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xix_xix_xpreheader_bbx_xnph7x_xix_xix_xi
      -- 	branch_block_stmt_2042/merge_stmt_3256__exit__
      -- 
    cp_elements(46) <= OrReduce(cp_elements(804) & cp_elements(826));
    -- CP-element group 47 place  bypass 
    -- predecessors 2024 
    -- successors 827 
    -- members (2) 
      -- 	branch_block_stmt_2042/assign_stmt_3278_to_assign_stmt_3283__entry__
      -- 	branch_block_stmt_2042/merge_stmt_3258__exit__
      -- 
    cp_elements(47) <= cp_elements(2024);
    -- CP-element group 48 merge  place  bypass 
    -- predecessors 837 841 
    -- successors 2045 
    -- members (2) 
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xix_xpreheader_bbx_xnphx_xix_xix_xi
      -- 	branch_block_stmt_2042/merge_stmt_3290__exit__
      -- 
    cp_elements(48) <= OrReduce(cp_elements(837) & cp_elements(841));
    -- CP-element group 49 place  bypass 
    -- predecessors 2067 
    -- successors 844 
    -- members (2) 
      -- 	branch_block_stmt_2042/assign_stmt_3312_to_assign_stmt_3323__entry__
      -- 	branch_block_stmt_2042/merge_stmt_3292__exit__
      -- 
    cp_elements(49) <= cp_elements(2067);
    -- CP-element group 50 branch  place  bypass 
    -- predecessors 858 
    -- successors 859 860 
    -- members (2) 
      -- 	branch_block_stmt_2042/if_stmt_3324__entry__
      -- 	branch_block_stmt_2042/assign_stmt_3312_to_assign_stmt_3323__exit__
      -- 
    cp_elements(50) <= cp_elements(858);
    -- CP-element group 51 merge  place  bypass 
    -- predecessors 859 2086 
    -- successors 2105 
    -- members (2) 
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xix_xloopexit_xx_x_crit_edgex_xix_xix_xi
      -- 	branch_block_stmt_2042/merge_stmt_3330__exit__
      -- 
    cp_elements(51) <= OrReduce(cp_elements(859) & cp_elements(2086));
    -- CP-element group 52 place  bypass 
    -- predecessors 2129 
    -- successors 866 
    -- members (2) 
      -- 	branch_block_stmt_2042/assign_stmt_3360_to_assign_stmt_3370__entry__
      -- 	branch_block_stmt_2042/merge_stmt_3341__exit__
      -- 
    cp_elements(52) <= cp_elements(2129);
    -- CP-element group 53 branch  place  bypass 
    -- predecessors 884 
    -- successors 885 886 
    -- members (2) 
      -- 	branch_block_stmt_2042/if_stmt_3371__entry__
      -- 	branch_block_stmt_2042/assign_stmt_3360_to_assign_stmt_3370__exit__
      -- 
    cp_elements(53) <= cp_elements(884);
    -- CP-element group 54 merge  fork  transition  place  bypass 
    -- predecessors 885 2135 
    -- successors 2139 2141 
    -- members (7) 
      -- 	branch_block_stmt_2042/merge_stmt_3377__exit__
      -- 	branch_block_stmt_2042/xx_xloopexitx_xix_xix_xix_xloopexit_xx_xloopexitx_xix_xix_xi
      -- 	branch_block_stmt_2042/xx_xloopexitx_xix_xix_xix_xloopexit_xx_xloopexitx_xix_xix_xi_PhiReq/phi_stmt_3385/phi_stmt_3385_sources/type_cast_3391/SplitProtocol/$entry
      -- 	branch_block_stmt_2042/xx_xloopexitx_xix_xix_xix_xloopexit_xx_xloopexitx_xix_xix_xi_PhiReq/phi_stmt_3385/phi_stmt_3385_sources/type_cast_3391/$entry
      -- 	branch_block_stmt_2042/xx_xloopexitx_xix_xix_xix_xloopexit_xx_xloopexitx_xix_xix_xi_PhiReq/phi_stmt_3385/phi_stmt_3385_sources/$entry
      -- 	branch_block_stmt_2042/xx_xloopexitx_xix_xix_xix_xloopexit_xx_xloopexitx_xix_xix_xi_PhiReq/phi_stmt_3385/$entry
      -- 	branch_block_stmt_2042/xx_xloopexitx_xix_xix_xix_xloopexit_xx_xloopexitx_xix_xix_xi_PhiReq/$entry
      -- 
    cp_elements(54) <= OrReduce(cp_elements(885) & cp_elements(2135));
    -- CP-element group 55 merge  place  bypass 
    -- predecessors 910 914 
    -- successors 2192 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xix_xpreheader_udiv32x_xexitx_xix_xi
      -- 	branch_block_stmt_2042/merge_stmt_3433__exit__
      -- 
    cp_elements(55) <= OrReduce(cp_elements(910) & cp_elements(914));
    -- CP-element group 56 place  bypass 
    -- predecessors 2214 
    -- successors 917 
    -- members (2) 
      -- 	branch_block_stmt_2042/assign_stmt_3455_to_assign_stmt_3486__entry__
      -- 	branch_block_stmt_2042/merge_stmt_3435__exit__
      -- 
    cp_elements(56) <= cp_elements(2214);
    -- CP-element group 57 branch  place  bypass 
    -- predecessors 943 
    -- successors 944 945 
    -- members (2) 
      -- 	branch_block_stmt_2042/if_stmt_3487__entry__
      -- 	branch_block_stmt_2042/assign_stmt_3455_to_assign_stmt_3486__exit__
      -- 
    cp_elements(57) <= cp_elements(943);
    -- CP-element group 58 merge  place  bypass 
    -- predecessors 944 2233 
    -- successors 951 
    -- members (2) 
      -- 	branch_block_stmt_2042/assign_stmt_3508_to_assign_stmt_3518__entry__
      -- 	branch_block_stmt_2042/merge_stmt_3493__exit__
      -- 
    cp_elements(58) <= OrReduce(cp_elements(944) & cp_elements(2233));
    -- CP-element group 59 place  bypass 
    -- predecessors 2290 
    -- successors 966 
    -- members (2) 
      -- 	branch_block_stmt_2042/assign_stmt_3539_to_assign_stmt_3565__entry__
      -- 	branch_block_stmt_2042/merge_stmt_3520__exit__
      -- 
    cp_elements(59) <= cp_elements(2290);
    -- CP-element group 60 merge  place  bypass 
    -- predecessors 1011 1017 
    -- successors 1018 
    -- members (2) 
      -- 	branch_block_stmt_2042/assign_stmt_3616__entry__
      -- 	branch_block_stmt_2042/merge_stmt_3610__exit__
      -- 
    cp_elements(60) <= OrReduce(cp_elements(1011) & cp_elements(1017));
    -- CP-element group 61 merge  fork  transition  place  bypass 
    -- predecessors 1023 1029 
    -- successors 2305 2307 
    -- members (7) 
      -- 	branch_block_stmt_2042/bb_57_bb_58
      -- 	branch_block_stmt_2042/merge_stmt_3623__exit__
      -- 	branch_block_stmt_2042/bb_57_bb_58_PhiReq/$entry
      -- 	branch_block_stmt_2042/bb_57_bb_58_PhiReq/phi_stmt_3626/$entry
      -- 	branch_block_stmt_2042/bb_57_bb_58_PhiReq/phi_stmt_3626/phi_stmt_3626_sources/$entry
      -- 	branch_block_stmt_2042/bb_57_bb_58_PhiReq/phi_stmt_3626/phi_stmt_3626_sources/type_cast_3629/$entry
      -- 	branch_block_stmt_2042/bb_57_bb_58_PhiReq/phi_stmt_3626/phi_stmt_3626_sources/type_cast_3629/SplitProtocol/$entry
      -- 
    cp_elements(61) <= OrReduce(cp_elements(1023) & cp_elements(1029));
    -- CP-element group 62 merge  place  bypass 
    -- predecessors 1043 1049 
    -- successors 1050 
    -- members (2) 
      -- 	branch_block_stmt_2042/merge_stmt_3660__exit__
      -- 	branch_block_stmt_2042/assign_stmt_3666__entry__
      -- 
    cp_elements(62) <= OrReduce(cp_elements(1043) & cp_elements(1049));
    -- CP-element group 63 merge  place  bypass 
    -- predecessors 1055 1061 
    -- successors 1062 
    -- members (2) 
      -- 	branch_block_stmt_2042/assign_stmt_3679__entry__
      -- 	branch_block_stmt_2042/merge_stmt_3673__exit__
      -- 
    cp_elements(63) <= OrReduce(cp_elements(1055) & cp_elements(1061));
    -- CP-element group 64 merge  place  bypass 
    -- predecessors 1067 2329 
    -- successors 1074 
    -- members (2) 
      -- 	branch_block_stmt_2042/assign_stmt_3701_to_assign_stmt_3719__entry__
      -- 	branch_block_stmt_2042/merge_stmt_3686__exit__
      -- 
    cp_elements(64) <= OrReduce(cp_elements(1067) & cp_elements(2329));
    -- CP-element group 65 place  bypass 
    -- predecessors 2372 
    -- successors 1088 
    -- members (2) 
      -- 	branch_block_stmt_2042/merge_stmt_3721__exit__
      -- 	branch_block_stmt_2042/assign_stmt_3741_to_assign_stmt_3747__entry__
      -- 
    cp_elements(65) <= cp_elements(2372);
    -- CP-element group 66 merge  place  bypass 
    -- predecessors 1096 1100 
    -- successors 2387 
    -- members (2) 
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xpreheader_bbx_xnphx_xix_xi
      -- 	branch_block_stmt_2042/merge_stmt_3754__exit__
      -- 
    cp_elements(66) <= OrReduce(cp_elements(1096) & cp_elements(1100));
    -- CP-element group 67 place  bypass 
    -- predecessors 2401 
    -- successors 1103 
    -- members (2) 
      -- 	branch_block_stmt_2042/merge_stmt_3756__exit__
      -- 	branch_block_stmt_2042/assign_stmt_3777_to_assign_stmt_3788__entry__
      -- 
    cp_elements(67) <= cp_elements(2401);
    -- CP-element group 68 branch  place  bypass 
    -- predecessors 1117 
    -- successors 1118 1119 
    -- members (2) 
      -- 	branch_block_stmt_2042/assign_stmt_3777_to_assign_stmt_3788__exit__
      -- 	branch_block_stmt_2042/if_stmt_3789__entry__
      -- 
    cp_elements(68) <= cp_elements(1117);
    -- CP-element group 69 merge  place  bypass 
    -- predecessors 1118 2420 
    -- successors 2431 
    -- members (2) 
      -- 	branch_block_stmt_2042/merge_stmt_3795__exit__
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xloopexit_xx_x_crit_edgex_xix_xi
      -- 
    cp_elements(69) <= OrReduce(cp_elements(1118) & cp_elements(2420));
    -- CP-element group 70 place  bypass 
    -- predecessors 2449 
    -- successors 1125 
    -- members (2) 
      -- 	branch_block_stmt_2042/merge_stmt_3806__exit__
      -- 	branch_block_stmt_2042/assign_stmt_3826_to_assign_stmt_3837__entry__
      -- 
    cp_elements(70) <= cp_elements(2449);
    -- CP-element group 71 branch  place  bypass 
    -- predecessors 1141 
    -- successors 1142 1143 
    -- members (2) 
      -- 	branch_block_stmt_2042/assign_stmt_3826_to_assign_stmt_3837__exit__
      -- 	branch_block_stmt_2042/if_stmt_3838__entry__
      -- 
    cp_elements(71) <= cp_elements(1141);
    -- CP-element group 72 merge  place  bypass 
    -- predecessors 1142 2455 
    -- successors 1149 
    -- members (2) 
      -- 	branch_block_stmt_2042/merge_stmt_3844__exit__
      -- 	branch_block_stmt_2042/assign_stmt_3855_to_assign_stmt_3898__entry__
      -- 
    cp_elements(72) <= OrReduce(cp_elements(1142) & cp_elements(2455));
    -- CP-element group 73 branch  place  bypass 
    -- predecessors 1181 
    -- successors 1182 1183 
    -- members (2) 
      -- 	branch_block_stmt_2042/assign_stmt_3855_to_assign_stmt_3898__exit__
      -- 	branch_block_stmt_2042/if_stmt_3899__entry__
      -- 
    cp_elements(73) <= cp_elements(1181);
    -- CP-element group 74 merge  place  bypass 
    -- predecessors 1182 1186 
    -- successors 2476 
    -- members (2) 
      -- 	branch_block_stmt_2042/merge_stmt_3905__exit__
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xpreheader_udiv32x_xexitx_xi
      -- 
    cp_elements(74) <= OrReduce(cp_elements(1182) & cp_elements(1186));
    -- CP-element group 75 place  bypass 
    -- predecessors 2498 
    -- successors 1189 
    -- members (2) 
      -- 	branch_block_stmt_2042/merge_stmt_3907__exit__
      -- 	branch_block_stmt_2042/assign_stmt_3927_to_assign_stmt_3958__entry__
      -- 
    cp_elements(75) <= cp_elements(2498);
    -- CP-element group 76 branch  place  bypass 
    -- predecessors 1215 
    -- successors 1216 1217 
    -- members (2) 
      -- 	branch_block_stmt_2042/assign_stmt_3927_to_assign_stmt_3958__exit__
      -- 	branch_block_stmt_2042/if_stmt_3959__entry__
      -- 
    cp_elements(76) <= cp_elements(1215);
    -- CP-element group 77 merge  place  bypass 
    -- predecessors 1216 2517 
    -- successors 1223 
    -- members (2) 
      -- 	branch_block_stmt_2042/merge_stmt_3965__exit__
      -- 	branch_block_stmt_2042/assign_stmt_3980_to_assign_stmt_3985__entry__
      -- 
    cp_elements(77) <= OrReduce(cp_elements(1216) & cp_elements(2517));
    -- CP-element group 78 place  bypass 
    -- predecessors 2574 
    -- successors 1233 
    -- members (2) 
      -- 	branch_block_stmt_2042/merge_stmt_3987__exit__
      -- 	branch_block_stmt_2042/assign_stmt_4006_to_assign_stmt_4032__entry__
      -- 
    cp_elements(78) <= cp_elements(2574);
    -- CP-element group 79 fork  transition  bypass 
    -- predecessors 2 
    -- successors 80 81 
    -- members (1) 
      -- 	branch_block_stmt_2042/assign_stmt_2069/$entry
      -- 
    cp_elements(79) <= cp_elements(2);
    -- CP-element group 80 transition  output  bypass 
    -- predecessors 79 
    -- successors 82 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_2069/RPIPE_in_data_2068_Sample/rr
      -- 	branch_block_stmt_2042/assign_stmt_2069/RPIPE_in_data_2068_Sample/$entry
      -- 	branch_block_stmt_2042/assign_stmt_2069/RPIPE_in_data_2068_sample_start_
      -- 
    cp_elements(80) <= cp_elements(79);
    rr_10614_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(80), ack => RPIPE_in_data_2068_inst_req_0); -- 
    -- CP-element group 81 transition  output  bypass 
    -- predecessors 79 
    -- successors 83 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_2069/RPIPE_in_data_2068_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_2069/RPIPE_in_data_2068_Update/$entry
      -- 	branch_block_stmt_2042/assign_stmt_2069/RPIPE_in_data_2068_Update/cr
      -- 
    cp_elements(81) <= cp_elements(79);
    cr_10619_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(81), ack => RPIPE_in_data_2068_inst_req_1); -- 
    -- CP-element group 82 transition  input  bypass 
    -- predecessors 80 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_2069/RPIPE_in_data_2068_Sample/$exit
      -- 	branch_block_stmt_2042/assign_stmt_2069/RPIPE_in_data_2068_Sample/ra
      -- 	branch_block_stmt_2042/assign_stmt_2069/RPIPE_in_data_2068_sample_completed_
      -- 
    ra_10615_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_in_data_2068_inst_ack_0, ack => cp_elements(82)); -- 
    -- CP-element group 83 transition  place  input  bypass 
    -- predecessors 81 
    -- successors 84 
    -- members (6) 
      -- 	branch_block_stmt_2042/assign_stmt_2069/RPIPE_in_data_2068_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2069/RPIPE_in_data_2068_Update/$exit
      -- 	branch_block_stmt_2042/assign_stmt_2069/RPIPE_in_data_2068_Update/ca
      -- 	branch_block_stmt_2042/assign_stmt_2069/$exit
      -- 	branch_block_stmt_2042/assign_stmt_2069__exit__
      -- 	branch_block_stmt_2042/assign_stmt_2072__entry__
      -- 
    ca_10620_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_in_data_2068_inst_ack_1, ack => cp_elements(83)); -- 
    -- CP-element group 84 fork  transition  bypass 
    -- predecessors 83 
    -- successors 85 86 
    -- members (1) 
      -- 	branch_block_stmt_2042/assign_stmt_2072/$entry
      -- 
    cp_elements(84) <= cp_elements(83);
    -- CP-element group 85 transition  output  bypass 
    -- predecessors 84 
    -- successors 87 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_2072/RPIPE_in_data_2071_Sample/$entry
      -- 	branch_block_stmt_2042/assign_stmt_2072/RPIPE_in_data_2071_Sample/rr
      -- 	branch_block_stmt_2042/assign_stmt_2072/RPIPE_in_data_2071_sample_start_
      -- 
    cp_elements(85) <= cp_elements(84);
    rr_10631_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(85), ack => RPIPE_in_data_2071_inst_req_0); -- 
    -- CP-element group 86 transition  output  bypass 
    -- predecessors 84 
    -- successors 88 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_2072/RPIPE_in_data_2071_Update/cr
      -- 	branch_block_stmt_2042/assign_stmt_2072/RPIPE_in_data_2071_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_2072/RPIPE_in_data_2071_Update/$entry
      -- 
    cp_elements(86) <= cp_elements(84);
    cr_10636_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(86), ack => RPIPE_in_data_2071_inst_req_1); -- 
    -- CP-element group 87 transition  input  bypass 
    -- predecessors 85 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_2072/RPIPE_in_data_2071_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2072/RPIPE_in_data_2071_Sample/$exit
      -- 	branch_block_stmt_2042/assign_stmt_2072/RPIPE_in_data_2071_Sample/ra
      -- 
    ra_10632_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_in_data_2071_inst_ack_0, ack => cp_elements(87)); -- 
    -- CP-element group 88 transition  place  input  bypass 
    -- predecessors 86 
    -- successors 89 
    -- members (6) 
      -- 	branch_block_stmt_2042/assign_stmt_2072/RPIPE_in_data_2071_Update/$exit
      -- 	branch_block_stmt_2042/assign_stmt_2072/RPIPE_in_data_2071_Update/ca
      -- 	branch_block_stmt_2042/assign_stmt_2072/RPIPE_in_data_2071_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2072/$exit
      -- 	branch_block_stmt_2042/assign_stmt_2072__exit__
      -- 	branch_block_stmt_2042/assign_stmt_2075__entry__
      -- 
    ca_10637_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_in_data_2071_inst_ack_1, ack => cp_elements(88)); -- 
    -- CP-element group 89 fork  transition  bypass 
    -- predecessors 88 
    -- successors 90 91 
    -- members (1) 
      -- 	branch_block_stmt_2042/assign_stmt_2075/$entry
      -- 
    cp_elements(89) <= cp_elements(88);
    -- CP-element group 90 transition  output  bypass 
    -- predecessors 89 
    -- successors 92 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_2075/RPIPE_in_data_2074_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_2075/RPIPE_in_data_2074_Sample/$entry
      -- 	branch_block_stmt_2042/assign_stmt_2075/RPIPE_in_data_2074_Sample/rr
      -- 
    cp_elements(90) <= cp_elements(89);
    rr_10648_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(90), ack => RPIPE_in_data_2074_inst_req_0); -- 
    -- CP-element group 91 transition  output  bypass 
    -- predecessors 89 
    -- successors 93 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_2075/RPIPE_in_data_2074_Update/cr
      -- 	branch_block_stmt_2042/assign_stmt_2075/RPIPE_in_data_2074_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_2075/RPIPE_in_data_2074_Update/$entry
      -- 
    cp_elements(91) <= cp_elements(89);
    cr_10653_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(91), ack => RPIPE_in_data_2074_inst_req_1); -- 
    -- CP-element group 92 transition  input  bypass 
    -- predecessors 90 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_2075/RPIPE_in_data_2074_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2075/RPIPE_in_data_2074_Sample/$exit
      -- 	branch_block_stmt_2042/assign_stmt_2075/RPIPE_in_data_2074_Sample/ra
      -- 
    ra_10649_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_in_data_2074_inst_ack_0, ack => cp_elements(92)); -- 
    -- CP-element group 93 transition  place  input  bypass 
    -- predecessors 91 
    -- successors 94 
    -- members (6) 
      -- 	branch_block_stmt_2042/assign_stmt_2075/RPIPE_in_data_2074_Update/$exit
      -- 	branch_block_stmt_2042/assign_stmt_2075/RPIPE_in_data_2074_Update/ca
      -- 	branch_block_stmt_2042/assign_stmt_2075/$exit
      -- 	branch_block_stmt_2042/assign_stmt_2075/RPIPE_in_data_2074_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2075__exit__
      -- 	branch_block_stmt_2042/assign_stmt_2078__entry__
      -- 
    ca_10654_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_in_data_2074_inst_ack_1, ack => cp_elements(93)); -- 
    -- CP-element group 94 fork  transition  bypass 
    -- predecessors 93 
    -- successors 95 96 
    -- members (1) 
      -- 	branch_block_stmt_2042/assign_stmt_2078/$entry
      -- 
    cp_elements(94) <= cp_elements(93);
    -- CP-element group 95 transition  output  bypass 
    -- predecessors 94 
    -- successors 97 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_2078/RPIPE_in_data_2077_Sample/rr
      -- 	branch_block_stmt_2042/assign_stmt_2078/RPIPE_in_data_2077_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_2078/RPIPE_in_data_2077_Sample/$entry
      -- 
    cp_elements(95) <= cp_elements(94);
    rr_10665_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(95), ack => RPIPE_in_data_2077_inst_req_0); -- 
    -- CP-element group 96 transition  output  bypass 
    -- predecessors 94 
    -- successors 98 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_2078/RPIPE_in_data_2077_Update/$entry
      -- 	branch_block_stmt_2042/assign_stmt_2078/RPIPE_in_data_2077_Update/cr
      -- 	branch_block_stmt_2042/assign_stmt_2078/RPIPE_in_data_2077_update_start_
      -- 
    cp_elements(96) <= cp_elements(94);
    cr_10670_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(96), ack => RPIPE_in_data_2077_inst_req_1); -- 
    -- CP-element group 97 transition  input  bypass 
    -- predecessors 95 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_2078/RPIPE_in_data_2077_Sample/$exit
      -- 	branch_block_stmt_2042/assign_stmt_2078/RPIPE_in_data_2077_Sample/ra
      -- 	branch_block_stmt_2042/assign_stmt_2078/RPIPE_in_data_2077_sample_completed_
      -- 
    ra_10666_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_in_data_2077_inst_ack_0, ack => cp_elements(97)); -- 
    -- CP-element group 98 transition  place  input  bypass 
    -- predecessors 96 
    -- successors 99 
    -- members (6) 
      -- 	branch_block_stmt_2042/assign_stmt_2078/RPIPE_in_data_2077_Update/ca
      -- 	branch_block_stmt_2042/assign_stmt_2078/RPIPE_in_data_2077_Update/$exit
      -- 	branch_block_stmt_2042/assign_stmt_2078/$exit
      -- 	branch_block_stmt_2042/assign_stmt_2078/RPIPE_in_data_2077_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2078__exit__
      -- 	branch_block_stmt_2042/assign_stmt_2083_to_assign_stmt_2111__entry__
      -- 
    ca_10671_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_in_data_2077_inst_ack_1, ack => cp_elements(98)); -- 
    -- CP-element group 99 fork  transition  bypass 
    -- predecessors 98 
    -- successors 101 102 103 106 110 111 114 117 120 
    -- members (1) 
      -- 	branch_block_stmt_2042/assign_stmt_2083_to_assign_stmt_2111/$entry
      -- 
    cp_elements(99) <= cp_elements(98);
    -- CP-element group 100 join  transition  output  bypass 
    -- predecessors 102 103 
    -- successors 104 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_2083_to_assign_stmt_2111/SUB_f32_f32_2082_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_2083_to_assign_stmt_2111/SUB_f32_f32_2082_Sample/rr
      -- 	branch_block_stmt_2042/assign_stmt_2083_to_assign_stmt_2111/SUB_f32_f32_2082_Sample/$entry
      -- 
    cp_element_group_100: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 20) := "cp_element_group_100"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(102) & cp_elements(103);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(100), clk => clk, reset => reset); --
    end block;
    rr_10690_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(100), ack => SUB_f32_f32_2082_inst_req_0); -- 
    -- CP-element group 101 transition  output  bypass 
    -- predecessors 99 
    -- successors 105 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_2083_to_assign_stmt_2111/SUB_f32_f32_2082_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_2083_to_assign_stmt_2111/SUB_f32_f32_2082_Update/$entry
      -- 	branch_block_stmt_2042/assign_stmt_2083_to_assign_stmt_2111/SUB_f32_f32_2082_Update/cr
      -- 
    cp_elements(101) <= cp_elements(99);
    cr_10695_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(101), ack => SUB_f32_f32_2082_inst_req_1); -- 
    -- CP-element group 102 transition  bypass 
    -- predecessors 99 
    -- successors 100 
    -- members (4) 
      -- 	branch_block_stmt_2042/assign_stmt_2083_to_assign_stmt_2111/R_iNsTr_8_2080_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_2083_to_assign_stmt_2111/R_iNsTr_8_2080_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2083_to_assign_stmt_2111/R_iNsTr_8_2080_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_2083_to_assign_stmt_2111/R_iNsTr_8_2080_update_completed_
      -- 
    cp_elements(102) <= cp_elements(99);
    -- CP-element group 103 transition  bypass 
    -- predecessors 99 
    -- successors 100 
    -- members (4) 
      -- 	branch_block_stmt_2042/assign_stmt_2083_to_assign_stmt_2111/R_iNsTr_6_2081_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_2083_to_assign_stmt_2111/R_iNsTr_6_2081_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2083_to_assign_stmt_2111/R_iNsTr_6_2081_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_2083_to_assign_stmt_2111/R_iNsTr_6_2081_update_completed_
      -- 
    cp_elements(103) <= cp_elements(99);
    -- CP-element group 104 transition  input  bypass 
    -- predecessors 100 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_2083_to_assign_stmt_2111/SUB_f32_f32_2082_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2083_to_assign_stmt_2111/SUB_f32_f32_2082_Sample/ra
      -- 	branch_block_stmt_2042/assign_stmt_2083_to_assign_stmt_2111/SUB_f32_f32_2082_Sample/$exit
      -- 
    ra_10691_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => SUB_f32_f32_2082_inst_ack_0, ack => cp_elements(104)); -- 
    -- CP-element group 105 transition  input  output  bypass 
    -- predecessors 101 
    -- successors 107 
    -- members (10) 
      -- 	branch_block_stmt_2042/assign_stmt_2083_to_assign_stmt_2111/MUL_f32_f32_2088_Sample/$entry
      -- 	branch_block_stmt_2042/assign_stmt_2083_to_assign_stmt_2111/MUL_f32_f32_2088_Sample/rr
      -- 	branch_block_stmt_2042/assign_stmt_2083_to_assign_stmt_2111/MUL_f32_f32_2088_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_2083_to_assign_stmt_2111/R_iNsTr_9_2085_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_2083_to_assign_stmt_2111/R_iNsTr_9_2085_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2083_to_assign_stmt_2111/R_iNsTr_9_2085_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_2083_to_assign_stmt_2111/R_iNsTr_9_2085_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2083_to_assign_stmt_2111/SUB_f32_f32_2082_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2083_to_assign_stmt_2111/SUB_f32_f32_2082_Update/$exit
      -- 	branch_block_stmt_2042/assign_stmt_2083_to_assign_stmt_2111/SUB_f32_f32_2082_Update/ca
      -- 
    ca_10696_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => SUB_f32_f32_2082_inst_ack_1, ack => cp_elements(105)); -- 
    rr_10708_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(105), ack => MUL_f32_f32_2088_inst_req_0); -- 
    -- CP-element group 106 transition  output  bypass 
    -- predecessors 99 
    -- successors 108 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_2083_to_assign_stmt_2111/MUL_f32_f32_2088_Update/cr
      -- 	branch_block_stmt_2042/assign_stmt_2083_to_assign_stmt_2111/MUL_f32_f32_2088_Update/$entry
      -- 	branch_block_stmt_2042/assign_stmt_2083_to_assign_stmt_2111/MUL_f32_f32_2088_update_start_
      -- 
    cp_elements(106) <= cp_elements(99);
    cr_10713_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(106), ack => MUL_f32_f32_2088_inst_req_1); -- 
    -- CP-element group 107 transition  input  bypass 
    -- predecessors 105 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_2083_to_assign_stmt_2111/MUL_f32_f32_2088_Sample/$exit
      -- 	branch_block_stmt_2042/assign_stmt_2083_to_assign_stmt_2111/MUL_f32_f32_2088_Sample/ra
      -- 	branch_block_stmt_2042/assign_stmt_2083_to_assign_stmt_2111/MUL_f32_f32_2088_sample_completed_
      -- 
    ra_10709_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => MUL_f32_f32_2088_inst_ack_0, ack => cp_elements(107)); -- 
    -- CP-element group 108 transition  input  bypass 
    -- predecessors 106 
    -- successors 109 
    -- members (7) 
      -- 	branch_block_stmt_2042/assign_stmt_2083_to_assign_stmt_2111/R_iNsTr_10_2091_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_2083_to_assign_stmt_2111/R_iNsTr_10_2091_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2083_to_assign_stmt_2111/R_iNsTr_10_2091_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_2083_to_assign_stmt_2111/R_iNsTr_10_2091_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2083_to_assign_stmt_2111/MUL_f32_f32_2088_Update/$exit
      -- 	branch_block_stmt_2042/assign_stmt_2083_to_assign_stmt_2111/MUL_f32_f32_2088_Update/ca
      -- 	branch_block_stmt_2042/assign_stmt_2083_to_assign_stmt_2111/MUL_f32_f32_2088_update_completed_
      -- 
    ca_10714_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => MUL_f32_f32_2088_inst_ack_1, ack => cp_elements(108)); -- 
    -- CP-element group 109 join  transition  output  bypass 
    -- predecessors 108 111 
    -- successors 112 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_2083_to_assign_stmt_2111/ADD_f32_f32_2093_Sample/$entry
      -- 	branch_block_stmt_2042/assign_stmt_2083_to_assign_stmt_2111/ADD_f32_f32_2093_Sample/rr
      -- 	branch_block_stmt_2042/assign_stmt_2083_to_assign_stmt_2111/ADD_f32_f32_2093_sample_start_
      -- 
    cp_element_group_109: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 20) := "cp_element_group_109"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(108) & cp_elements(111);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(109), clk => clk, reset => reset); --
    end block;
    rr_10730_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(109), ack => ADD_f32_f32_2093_inst_req_0); -- 
    -- CP-element group 110 transition  output  bypass 
    -- predecessors 99 
    -- successors 113 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_2083_to_assign_stmt_2111/ADD_f32_f32_2093_Update/$entry
      -- 	branch_block_stmt_2042/assign_stmt_2083_to_assign_stmt_2111/ADD_f32_f32_2093_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_2083_to_assign_stmt_2111/ADD_f32_f32_2093_Update/cr
      -- 
    cp_elements(110) <= cp_elements(99);
    cr_10735_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(110), ack => ADD_f32_f32_2093_inst_req_1); -- 
    -- CP-element group 111 transition  bypass 
    -- predecessors 99 
    -- successors 109 
    -- members (4) 
      -- 	branch_block_stmt_2042/assign_stmt_2083_to_assign_stmt_2111/R_int_speed_errx_x0_2092_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_2083_to_assign_stmt_2111/R_int_speed_errx_x0_2092_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2083_to_assign_stmt_2111/R_int_speed_errx_x0_2092_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_2083_to_assign_stmt_2111/R_int_speed_errx_x0_2092_sample_completed_
      -- 
    cp_elements(111) <= cp_elements(99);
    -- CP-element group 112 transition  input  bypass 
    -- predecessors 109 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_2083_to_assign_stmt_2111/ADD_f32_f32_2093_Sample/$exit
      -- 	branch_block_stmt_2042/assign_stmt_2083_to_assign_stmt_2111/ADD_f32_f32_2093_Sample/ra
      -- 	branch_block_stmt_2042/assign_stmt_2083_to_assign_stmt_2111/ADD_f32_f32_2093_sample_completed_
      -- 
    ra_10731_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_f32_f32_2093_inst_ack_0, ack => cp_elements(112)); -- 
    -- CP-element group 113 transition  input  output  bypass 
    -- predecessors 110 
    -- successors 115 
    -- members (10) 
      -- 	branch_block_stmt_2042/assign_stmt_2083_to_assign_stmt_2111/MUL_f32_f32_2099_Sample/rr
      -- 	branch_block_stmt_2042/assign_stmt_2083_to_assign_stmt_2111/ADD_f32_f32_2093_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2083_to_assign_stmt_2111/R_iNsTr_11_2096_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2083_to_assign_stmt_2111/MUL_f32_f32_2099_Sample/$entry
      -- 	branch_block_stmt_2042/assign_stmt_2083_to_assign_stmt_2111/MUL_f32_f32_2099_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_2083_to_assign_stmt_2111/R_iNsTr_11_2096_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_2083_to_assign_stmt_2111/R_iNsTr_11_2096_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2083_to_assign_stmt_2111/R_iNsTr_11_2096_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_2083_to_assign_stmt_2111/ADD_f32_f32_2093_Update/$exit
      -- 	branch_block_stmt_2042/assign_stmt_2083_to_assign_stmt_2111/ADD_f32_f32_2093_Update/ca
      -- 
    ca_10736_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_f32_f32_2093_inst_ack_1, ack => cp_elements(113)); -- 
    rr_10748_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(113), ack => MUL_f32_f32_2099_inst_req_0); -- 
    -- CP-element group 114 transition  output  bypass 
    -- predecessors 99 
    -- successors 116 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_2083_to_assign_stmt_2111/MUL_f32_f32_2099_Update/$entry
      -- 	branch_block_stmt_2042/assign_stmt_2083_to_assign_stmt_2111/MUL_f32_f32_2099_Update/cr
      -- 	branch_block_stmt_2042/assign_stmt_2083_to_assign_stmt_2111/MUL_f32_f32_2099_update_start_
      -- 
    cp_elements(114) <= cp_elements(99);
    cr_10753_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(114), ack => MUL_f32_f32_2099_inst_req_1); -- 
    -- CP-element group 115 transition  input  bypass 
    -- predecessors 113 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_2083_to_assign_stmt_2111/MUL_f32_f32_2099_Sample/$exit
      -- 	branch_block_stmt_2042/assign_stmt_2083_to_assign_stmt_2111/MUL_f32_f32_2099_Sample/ra
      -- 	branch_block_stmt_2042/assign_stmt_2083_to_assign_stmt_2111/MUL_f32_f32_2099_sample_completed_
      -- 
    ra_10749_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => MUL_f32_f32_2099_inst_ack_0, ack => cp_elements(115)); -- 
    -- CP-element group 116 transition  input  output  bypass 
    -- predecessors 114 
    -- successors 118 
    -- members (10) 
      -- 	branch_block_stmt_2042/assign_stmt_2083_to_assign_stmt_2111/type_cast_2104_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_2083_to_assign_stmt_2111/R_iNsTr_12_2103_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_2083_to_assign_stmt_2111/R_iNsTr_12_2103_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2083_to_assign_stmt_2111/R_iNsTr_12_2103_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_2083_to_assign_stmt_2111/MUL_f32_f32_2099_Update/$exit
      -- 	branch_block_stmt_2042/assign_stmt_2083_to_assign_stmt_2111/MUL_f32_f32_2099_Update/ca
      -- 	branch_block_stmt_2042/assign_stmt_2083_to_assign_stmt_2111/type_cast_2104_Sample/$entry
      -- 	branch_block_stmt_2042/assign_stmt_2083_to_assign_stmt_2111/type_cast_2104_Sample/rr
      -- 	branch_block_stmt_2042/assign_stmt_2083_to_assign_stmt_2111/MUL_f32_f32_2099_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2083_to_assign_stmt_2111/R_iNsTr_12_2103_update_completed_
      -- 
    ca_10754_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => MUL_f32_f32_2099_inst_ack_1, ack => cp_elements(116)); -- 
    rr_10766_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(116), ack => type_cast_2104_inst_req_0); -- 
    -- CP-element group 117 transition  output  bypass 
    -- predecessors 99 
    -- successors 119 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_2083_to_assign_stmt_2111/type_cast_2104_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_2083_to_assign_stmt_2111/type_cast_2104_Update/$entry
      -- 	branch_block_stmt_2042/assign_stmt_2083_to_assign_stmt_2111/type_cast_2104_Update/cr
      -- 
    cp_elements(117) <= cp_elements(99);
    cr_10771_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(117), ack => type_cast_2104_inst_req_1); -- 
    -- CP-element group 118 transition  input  bypass 
    -- predecessors 116 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_2083_to_assign_stmt_2111/type_cast_2104_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2083_to_assign_stmt_2111/type_cast_2104_Sample/$exit
      -- 	branch_block_stmt_2042/assign_stmt_2083_to_assign_stmt_2111/type_cast_2104_Sample/ra
      -- 
    ra_10767_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2104_inst_ack_0, ack => cp_elements(118)); -- 
    -- CP-element group 119 transition  input  output  bypass 
    -- predecessors 117 
    -- successors 121 
    -- members (10) 
      -- 	branch_block_stmt_2042/assign_stmt_2083_to_assign_stmt_2111/R_iNsTr_13_2107_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2083_to_assign_stmt_2111/type_cast_2104_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2083_to_assign_stmt_2111/SLT_f64_u1_2110_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_2083_to_assign_stmt_2111/R_iNsTr_13_2107_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_2083_to_assign_stmt_2111/R_iNsTr_13_2107_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2083_to_assign_stmt_2111/R_iNsTr_13_2107_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_2083_to_assign_stmt_2111/type_cast_2104_Update/$exit
      -- 	branch_block_stmt_2042/assign_stmt_2083_to_assign_stmt_2111/type_cast_2104_Update/ca
      -- 	branch_block_stmt_2042/assign_stmt_2083_to_assign_stmt_2111/SLT_f64_u1_2110_Sample/$entry
      -- 	branch_block_stmt_2042/assign_stmt_2083_to_assign_stmt_2111/SLT_f64_u1_2110_Sample/rr
      -- 
    ca_10772_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2104_inst_ack_1, ack => cp_elements(119)); -- 
    rr_10784_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(119), ack => SLT_f64_u1_2110_inst_req_0); -- 
    -- CP-element group 120 transition  output  bypass 
    -- predecessors 99 
    -- successors 122 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_2083_to_assign_stmt_2111/SLT_f64_u1_2110_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_2083_to_assign_stmt_2111/SLT_f64_u1_2110_Update/$entry
      -- 	branch_block_stmt_2042/assign_stmt_2083_to_assign_stmt_2111/SLT_f64_u1_2110_Update/cr
      -- 
    cp_elements(120) <= cp_elements(99);
    cr_10789_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(120), ack => SLT_f64_u1_2110_inst_req_1); -- 
    -- CP-element group 121 transition  input  bypass 
    -- predecessors 119 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_2083_to_assign_stmt_2111/SLT_f64_u1_2110_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2083_to_assign_stmt_2111/SLT_f64_u1_2110_Sample/$exit
      -- 	branch_block_stmt_2042/assign_stmt_2083_to_assign_stmt_2111/SLT_f64_u1_2110_Sample/ra
      -- 
    ra_10785_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => SLT_f64_u1_2110_inst_ack_0, ack => cp_elements(121)); -- 
    -- CP-element group 122 branch  transition  place  input  bypass 
    -- predecessors 120 
    -- successors 123 124 
    -- members (6) 
      -- 	branch_block_stmt_2042/assign_stmt_2083_to_assign_stmt_2111/SLT_f64_u1_2110_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2083_to_assign_stmt_2111/$exit
      -- 	branch_block_stmt_2042/assign_stmt_2083_to_assign_stmt_2111/SLT_f64_u1_2110_Update/ca
      -- 	branch_block_stmt_2042/assign_stmt_2083_to_assign_stmt_2111/SLT_f64_u1_2110_Update/$exit
      -- 	branch_block_stmt_2042/assign_stmt_2083_to_assign_stmt_2111__exit__
      -- 	branch_block_stmt_2042/if_stmt_2112__entry__
      -- 
    ca_10790_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => SLT_f64_u1_2110_inst_ack_1, ack => cp_elements(122)); -- 
    -- CP-element group 123 transition  place  dead  bypass 
    -- predecessors 122 
    -- successors 3 
    -- members (8) 
      -- 	branch_block_stmt_2042/if_stmt_2112_dead_link/$entry
      -- 	branch_block_stmt_2042/if_stmt_2112_dead_link/$exit
      -- 	branch_block_stmt_2042/if_stmt_2112_dead_link/dead_transition
      -- 	branch_block_stmt_2042/if_stmt_2112__exit__
      -- 	branch_block_stmt_2042/merge_stmt_2118__entry__
      -- 	branch_block_stmt_2042/merge_stmt_2118_dead_link/$entry
      -- 	branch_block_stmt_2042/merge_stmt_2118_dead_link/$exit
      -- 	branch_block_stmt_2042/merge_stmt_2118_dead_link/dead_transition
      -- 
    cp_elements(123) <= false;
    -- CP-element group 124 transition  output  bypass 
    -- predecessors 122 
    -- successors 125 
    -- members (3) 
      -- 	branch_block_stmt_2042/if_stmt_2112_eval_test/$entry
      -- 	branch_block_stmt_2042/if_stmt_2112_eval_test/$exit
      -- 	branch_block_stmt_2042/if_stmt_2112_eval_test/branch_req
      -- 
    cp_elements(124) <= cp_elements(122);
    branch_req_10798_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(124), ack => if_stmt_2112_branch_req_0); -- 
    -- CP-element group 125 branch  place  bypass 
    -- predecessors 124 
    -- successors 126 128 
    -- members (1) 
      -- 	branch_block_stmt_2042/R_iNsTr_14_2113_place
      -- 
    cp_elements(125) <= cp_elements(124);
    -- CP-element group 126 transition  bypass 
    -- predecessors 125 
    -- successors 127 
    -- members (1) 
      -- 	branch_block_stmt_2042/if_stmt_2112_if_link/$entry
      -- 
    cp_elements(126) <= cp_elements(125);
    -- CP-element group 127 fork  transition  place  input  bypass 
    -- predecessors 126 
    -- successors 1317 1318 
    -- members (8) 
      -- 	branch_block_stmt_2042/bb_1_bb_4
      -- 	branch_block_stmt_2042/if_stmt_2112_if_link/$exit
      -- 	branch_block_stmt_2042/if_stmt_2112_if_link/if_choice_transition
      -- 	branch_block_stmt_2042/bb_1_bb_4_PhiReq/$entry
      -- 	branch_block_stmt_2042/bb_1_bb_4_PhiReq/phi_stmt_2134/$entry
      -- 	branch_block_stmt_2042/bb_1_bb_4_PhiReq/phi_stmt_2134/phi_stmt_2134_sources/$entry
      -- 	branch_block_stmt_2042/bb_1_bb_4_PhiReq/phi_stmt_2134/phi_stmt_2134_sources/type_cast_2137/$entry
      -- 	branch_block_stmt_2042/bb_1_bb_4_PhiReq/phi_stmt_2134/phi_stmt_2134_sources/type_cast_2137/SplitProtocol/$entry
      -- 
    if_choice_transition_10803_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2112_branch_ack_1, ack => cp_elements(127)); -- 
    -- CP-element group 128 transition  bypass 
    -- predecessors 125 
    -- successors 129 
    -- members (1) 
      -- 	branch_block_stmt_2042/if_stmt_2112_else_link/$entry
      -- 
    cp_elements(128) <= cp_elements(125);
    -- CP-element group 129 transition  place  input  bypass 
    -- predecessors 128 
    -- successors 3 
    -- members (9) 
      -- 	branch_block_stmt_2042/bb_1_bb_2
      -- 	branch_block_stmt_2042/if_stmt_2112_else_link/$exit
      -- 	branch_block_stmt_2042/if_stmt_2112_else_link/else_choice_transition
      -- 	branch_block_stmt_2042/merge_stmt_2118_PhiReqMerge
      -- 	branch_block_stmt_2042/bb_1_bb_2_PhiReq/$entry
      -- 	branch_block_stmt_2042/bb_1_bb_2_PhiReq/$exit
      -- 	branch_block_stmt_2042/merge_stmt_2118_PhiAck/$entry
      -- 	branch_block_stmt_2042/merge_stmt_2118_PhiAck/$exit
      -- 	branch_block_stmt_2042/merge_stmt_2118_PhiAck/dummy
      -- 
    else_choice_transition_10807_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2112_branch_ack_0, ack => cp_elements(129)); -- 
    -- CP-element group 130 fork  transition  bypass 
    -- predecessors 3 
    -- successors 131 132 
    -- members (1) 
      -- 	branch_block_stmt_2042/assign_stmt_2124/$entry
      -- 
    cp_elements(130) <= cp_elements(3);
    -- CP-element group 131 transition  output  bypass 
    -- predecessors 130 
    -- successors 134 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_2124/SGT_f64_u1_2123_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_2124/SGT_f64_u1_2123_Update/$entry
      -- 	branch_block_stmt_2042/assign_stmt_2124/SGT_f64_u1_2123_Update/cr
      -- 
    cp_elements(131) <= cp_elements(130);
    cr_10829_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(131), ack => SGT_f64_u1_2123_inst_req_1); -- 
    -- CP-element group 132 transition  output  bypass 
    -- predecessors 130 
    -- successors 133 
    -- members (7) 
      -- 	branch_block_stmt_2042/assign_stmt_2124/SGT_f64_u1_2123_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_2124/R_iNsTr_13_2120_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_2124/R_iNsTr_13_2120_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2124/R_iNsTr_13_2120_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_2124/R_iNsTr_13_2120_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2124/SGT_f64_u1_2123_Sample/$entry
      -- 	branch_block_stmt_2042/assign_stmt_2124/SGT_f64_u1_2123_Sample/rr
      -- 
    cp_elements(132) <= cp_elements(130);
    rr_10824_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(132), ack => SGT_f64_u1_2123_inst_req_0); -- 
    -- CP-element group 133 transition  input  bypass 
    -- predecessors 132 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_2124/SGT_f64_u1_2123_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2124/SGT_f64_u1_2123_Sample/$exit
      -- 	branch_block_stmt_2042/assign_stmt_2124/SGT_f64_u1_2123_Sample/ra
      -- 
    ra_10825_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => SGT_f64_u1_2123_inst_ack_0, ack => cp_elements(133)); -- 
    -- CP-element group 134 branch  transition  place  input  bypass 
    -- predecessors 131 
    -- successors 135 136 
    -- members (6) 
      -- 	branch_block_stmt_2042/assign_stmt_2124__exit__
      -- 	branch_block_stmt_2042/if_stmt_2125__entry__
      -- 	branch_block_stmt_2042/assign_stmt_2124/$exit
      -- 	branch_block_stmt_2042/assign_stmt_2124/SGT_f64_u1_2123_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2124/SGT_f64_u1_2123_Update/$exit
      -- 	branch_block_stmt_2042/assign_stmt_2124/SGT_f64_u1_2123_Update/ca
      -- 
    ca_10830_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => SGT_f64_u1_2123_inst_ack_1, ack => cp_elements(134)); -- 
    -- CP-element group 135 transition  place  dead  bypass 
    -- predecessors 134 
    -- successors 4 
    -- members (8) 
      -- 	branch_block_stmt_2042/if_stmt_2125__exit__
      -- 	branch_block_stmt_2042/merge_stmt_2131__entry__
      -- 	branch_block_stmt_2042/if_stmt_2125_dead_link/$entry
      -- 	branch_block_stmt_2042/if_stmt_2125_dead_link/$exit
      -- 	branch_block_stmt_2042/if_stmt_2125_dead_link/dead_transition
      -- 	branch_block_stmt_2042/merge_stmt_2131_dead_link/$entry
      -- 	branch_block_stmt_2042/merge_stmt_2131_dead_link/$exit
      -- 	branch_block_stmt_2042/merge_stmt_2131_dead_link/dead_transition
      -- 
    cp_elements(135) <= false;
    -- CP-element group 136 transition  output  bypass 
    -- predecessors 134 
    -- successors 137 
    -- members (3) 
      -- 	branch_block_stmt_2042/if_stmt_2125_eval_test/$entry
      -- 	branch_block_stmt_2042/if_stmt_2125_eval_test/$exit
      -- 	branch_block_stmt_2042/if_stmt_2125_eval_test/branch_req
      -- 
    cp_elements(136) <= cp_elements(134);
    branch_req_10838_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(136), ack => if_stmt_2125_branch_req_0); -- 
    -- CP-element group 137 branch  place  bypass 
    -- predecessors 136 
    -- successors 138 140 
    -- members (1) 
      -- 	branch_block_stmt_2042/R_iNsTr_20_2126_place
      -- 
    cp_elements(137) <= cp_elements(136);
    -- CP-element group 138 transition  bypass 
    -- predecessors 137 
    -- successors 139 
    -- members (1) 
      -- 	branch_block_stmt_2042/if_stmt_2125_if_link/$entry
      -- 
    cp_elements(138) <= cp_elements(137);
    -- CP-element group 139 fork  transition  place  input  bypass 
    -- predecessors 138 
    -- successors 1320 1321 
    -- members (8) 
      -- 	branch_block_stmt_2042/if_stmt_2125_if_link/$exit
      -- 	branch_block_stmt_2042/if_stmt_2125_if_link/if_choice_transition
      -- 	branch_block_stmt_2042/bb_2_bb_4
      -- 	branch_block_stmt_2042/bb_2_bb_4_PhiReq/$entry
      -- 	branch_block_stmt_2042/bb_2_bb_4_PhiReq/phi_stmt_2134/$entry
      -- 	branch_block_stmt_2042/bb_2_bb_4_PhiReq/phi_stmt_2134/phi_stmt_2134_sources/$entry
      -- 	branch_block_stmt_2042/bb_2_bb_4_PhiReq/phi_stmt_2134/phi_stmt_2134_sources/type_cast_2137/$entry
      -- 	branch_block_stmt_2042/bb_2_bb_4_PhiReq/phi_stmt_2134/phi_stmt_2134_sources/type_cast_2137/SplitProtocol/$entry
      -- 
    if_choice_transition_10843_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2125_branch_ack_1, ack => cp_elements(139)); -- 
    -- CP-element group 140 transition  bypass 
    -- predecessors 137 
    -- successors 141 
    -- members (1) 
      -- 	branch_block_stmt_2042/if_stmt_2125_else_link/$entry
      -- 
    cp_elements(140) <= cp_elements(137);
    -- CP-element group 141 transition  place  input  bypass 
    -- predecessors 140 
    -- successors 4 
    -- members (9) 
      -- 	branch_block_stmt_2042/if_stmt_2125_else_link/$exit
      -- 	branch_block_stmt_2042/if_stmt_2125_else_link/else_choice_transition
      -- 	branch_block_stmt_2042/bb_2_bb_3
      -- 	branch_block_stmt_2042/merge_stmt_2131_PhiReqMerge
      -- 	branch_block_stmt_2042/bb_2_bb_3_PhiReq/$entry
      -- 	branch_block_stmt_2042/bb_2_bb_3_PhiReq/$exit
      -- 	branch_block_stmt_2042/merge_stmt_2131_PhiAck/$entry
      -- 	branch_block_stmt_2042/merge_stmt_2131_PhiAck/$exit
      -- 	branch_block_stmt_2042/merge_stmt_2131_PhiAck/dummy
      -- 
    else_choice_transition_10847_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2125_branch_ack_0, ack => cp_elements(141)); -- 
    -- CP-element group 142 fork  transition  bypass 
    -- predecessors 1330 
    -- successors 143 144 148 149 152 
    -- members (1) 
      -- 	branch_block_stmt_2042/assign_stmt_2150_to_assign_stmt_2161/$entry
      -- 
    cp_elements(142) <= cp_elements(1330);
    -- CP-element group 143 transition  output  bypass 
    -- predecessors 142 
    -- successors 146 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_2150_to_assign_stmt_2161/MUL_f32_f32_2149_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_2150_to_assign_stmt_2161/MUL_f32_f32_2149_Update/$entry
      -- 	branch_block_stmt_2042/assign_stmt_2150_to_assign_stmt_2161/MUL_f32_f32_2149_Update/cr
      -- 
    cp_elements(143) <= cp_elements(142);
    cr_10869_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(143), ack => MUL_f32_f32_2149_inst_req_1); -- 
    -- CP-element group 144 transition  output  bypass 
    -- predecessors 142 
    -- successors 145 
    -- members (7) 
      -- 	branch_block_stmt_2042/assign_stmt_2150_to_assign_stmt_2161/MUL_f32_f32_2149_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_2150_to_assign_stmt_2161/R_iNsTr_9_2146_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_2150_to_assign_stmt_2161/R_iNsTr_9_2146_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2150_to_assign_stmt_2161/R_iNsTr_9_2146_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_2150_to_assign_stmt_2161/R_iNsTr_9_2146_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2150_to_assign_stmt_2161/MUL_f32_f32_2149_Sample/$entry
      -- 	branch_block_stmt_2042/assign_stmt_2150_to_assign_stmt_2161/MUL_f32_f32_2149_Sample/rr
      -- 
    cp_elements(144) <= cp_elements(142);
    rr_10864_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(144), ack => MUL_f32_f32_2149_inst_req_0); -- 
    -- CP-element group 145 transition  input  bypass 
    -- predecessors 144 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_2150_to_assign_stmt_2161/MUL_f32_f32_2149_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2150_to_assign_stmt_2161/MUL_f32_f32_2149_Sample/$exit
      -- 	branch_block_stmt_2042/assign_stmt_2150_to_assign_stmt_2161/MUL_f32_f32_2149_Sample/ra
      -- 
    ra_10865_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => MUL_f32_f32_2149_inst_ack_0, ack => cp_elements(145)); -- 
    -- CP-element group 146 transition  input  bypass 
    -- predecessors 143 
    -- successors 147 
    -- members (7) 
      -- 	branch_block_stmt_2042/assign_stmt_2150_to_assign_stmt_2161/MUL_f32_f32_2149_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2150_to_assign_stmt_2161/MUL_f32_f32_2149_Update/$exit
      -- 	branch_block_stmt_2042/assign_stmt_2150_to_assign_stmt_2161/MUL_f32_f32_2149_Update/ca
      -- 	branch_block_stmt_2042/assign_stmt_2150_to_assign_stmt_2161/R_iNsTr_16_2153_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_2150_to_assign_stmt_2161/R_iNsTr_16_2153_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2150_to_assign_stmt_2161/R_iNsTr_16_2153_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_2150_to_assign_stmt_2161/R_iNsTr_16_2153_update_completed_
      -- 
    ca_10870_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => MUL_f32_f32_2149_inst_ack_1, ack => cp_elements(146)); -- 
    -- CP-element group 147 join  transition  output  bypass 
    -- predecessors 146 149 
    -- successors 150 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_2150_to_assign_stmt_2161/ADD_f32_f32_2154_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_2150_to_assign_stmt_2161/ADD_f32_f32_2154_Sample/$entry
      -- 	branch_block_stmt_2042/assign_stmt_2150_to_assign_stmt_2161/ADD_f32_f32_2154_Sample/rr
      -- 
    cp_element_group_147: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 20) := "cp_element_group_147"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(146) & cp_elements(149);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(147), clk => clk, reset => reset); --
    end block;
    rr_10886_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(147), ack => ADD_f32_f32_2154_inst_req_0); -- 
    -- CP-element group 148 transition  output  bypass 
    -- predecessors 142 
    -- successors 151 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_2150_to_assign_stmt_2161/ADD_f32_f32_2154_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_2150_to_assign_stmt_2161/ADD_f32_f32_2154_Update/$entry
      -- 	branch_block_stmt_2042/assign_stmt_2150_to_assign_stmt_2161/ADD_f32_f32_2154_Update/cr
      -- 
    cp_elements(148) <= cp_elements(142);
    cr_10891_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(148), ack => ADD_f32_f32_2154_inst_req_1); -- 
    -- CP-element group 149 transition  bypass 
    -- predecessors 142 
    -- successors 147 
    -- members (4) 
      -- 	branch_block_stmt_2042/assign_stmt_2150_to_assign_stmt_2161/R_int_speed_errx_x1_2152_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_2150_to_assign_stmt_2161/R_int_speed_errx_x1_2152_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2150_to_assign_stmt_2161/R_int_speed_errx_x1_2152_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_2150_to_assign_stmt_2161/R_int_speed_errx_x1_2152_update_completed_
      -- 
    cp_elements(149) <= cp_elements(142);
    -- CP-element group 150 transition  input  bypass 
    -- predecessors 147 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_2150_to_assign_stmt_2161/ADD_f32_f32_2154_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2150_to_assign_stmt_2161/ADD_f32_f32_2154_Sample/$exit
      -- 	branch_block_stmt_2042/assign_stmt_2150_to_assign_stmt_2161/ADD_f32_f32_2154_Sample/ra
      -- 
    ra_10887_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_f32_f32_2154_inst_ack_0, ack => cp_elements(150)); -- 
    -- CP-element group 151 transition  input  output  bypass 
    -- predecessors 148 
    -- successors 153 
    -- members (10) 
      -- 	branch_block_stmt_2042/assign_stmt_2150_to_assign_stmt_2161/ADD_f32_f32_2154_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2150_to_assign_stmt_2161/ADD_f32_f32_2154_Update/$exit
      -- 	branch_block_stmt_2042/assign_stmt_2150_to_assign_stmt_2161/ADD_f32_f32_2154_Update/ca
      -- 	branch_block_stmt_2042/assign_stmt_2150_to_assign_stmt_2161/SLT_f32_u1_2160_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_2150_to_assign_stmt_2161/R_iNsTr_17_2157_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_2150_to_assign_stmt_2161/R_iNsTr_17_2157_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2150_to_assign_stmt_2161/R_iNsTr_17_2157_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_2150_to_assign_stmt_2161/R_iNsTr_17_2157_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2150_to_assign_stmt_2161/SLT_f32_u1_2160_Sample/$entry
      -- 	branch_block_stmt_2042/assign_stmt_2150_to_assign_stmt_2161/SLT_f32_u1_2160_Sample/rr
      -- 
    ca_10892_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_f32_f32_2154_inst_ack_1, ack => cp_elements(151)); -- 
    rr_10904_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(151), ack => SLT_f32_u1_2160_inst_req_0); -- 
    -- CP-element group 152 transition  output  bypass 
    -- predecessors 142 
    -- successors 154 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_2150_to_assign_stmt_2161/SLT_f32_u1_2160_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_2150_to_assign_stmt_2161/SLT_f32_u1_2160_Update/$entry
      -- 	branch_block_stmt_2042/assign_stmt_2150_to_assign_stmt_2161/SLT_f32_u1_2160_Update/cr
      -- 
    cp_elements(152) <= cp_elements(142);
    cr_10909_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(152), ack => SLT_f32_u1_2160_inst_req_1); -- 
    -- CP-element group 153 transition  input  bypass 
    -- predecessors 151 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_2150_to_assign_stmt_2161/SLT_f32_u1_2160_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2150_to_assign_stmt_2161/SLT_f32_u1_2160_Sample/$exit
      -- 	branch_block_stmt_2042/assign_stmt_2150_to_assign_stmt_2161/SLT_f32_u1_2160_Sample/ra
      -- 
    ra_10905_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => SLT_f32_u1_2160_inst_ack_0, ack => cp_elements(153)); -- 
    -- CP-element group 154 branch  transition  place  input  bypass 
    -- predecessors 152 
    -- successors 155 156 
    -- members (6) 
      -- 	branch_block_stmt_2042/assign_stmt_2150_to_assign_stmt_2161__exit__
      -- 	branch_block_stmt_2042/if_stmt_2162__entry__
      -- 	branch_block_stmt_2042/assign_stmt_2150_to_assign_stmt_2161/$exit
      -- 	branch_block_stmt_2042/assign_stmt_2150_to_assign_stmt_2161/SLT_f32_u1_2160_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2150_to_assign_stmt_2161/SLT_f32_u1_2160_Update/$exit
      -- 	branch_block_stmt_2042/assign_stmt_2150_to_assign_stmt_2161/SLT_f32_u1_2160_Update/ca
      -- 
    ca_10910_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => SLT_f32_u1_2160_inst_ack_1, ack => cp_elements(154)); -- 
    -- CP-element group 155 transition  place  dead  bypass 
    -- predecessors 154 
    -- successors 5 
    -- members (8) 
      -- 	branch_block_stmt_2042/if_stmt_2162__exit__
      -- 	branch_block_stmt_2042/merge_stmt_2168__entry__
      -- 	branch_block_stmt_2042/if_stmt_2162_dead_link/$entry
      -- 	branch_block_stmt_2042/if_stmt_2162_dead_link/$exit
      -- 	branch_block_stmt_2042/if_stmt_2162_dead_link/dead_transition
      -- 	branch_block_stmt_2042/merge_stmt_2168_dead_link/$entry
      -- 	branch_block_stmt_2042/merge_stmt_2168_dead_link/$exit
      -- 	branch_block_stmt_2042/merge_stmt_2168_dead_link/dead_transition
      -- 
    cp_elements(155) <= false;
    -- CP-element group 156 transition  output  bypass 
    -- predecessors 154 
    -- successors 157 
    -- members (3) 
      -- 	branch_block_stmt_2042/if_stmt_2162_eval_test/$entry
      -- 	branch_block_stmt_2042/if_stmt_2162_eval_test/$exit
      -- 	branch_block_stmt_2042/if_stmt_2162_eval_test/branch_req
      -- 
    cp_elements(156) <= cp_elements(154);
    branch_req_10918_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(156), ack => if_stmt_2162_branch_req_0); -- 
    -- CP-element group 157 branch  place  bypass 
    -- predecessors 156 
    -- successors 158 160 
    -- members (1) 
      -- 	branch_block_stmt_2042/R_iNsTr_18_2163_place
      -- 
    cp_elements(157) <= cp_elements(156);
    -- CP-element group 158 transition  bypass 
    -- predecessors 157 
    -- successors 159 
    -- members (1) 
      -- 	branch_block_stmt_2042/if_stmt_2162_if_link/$entry
      -- 
    cp_elements(158) <= cp_elements(157);
    -- CP-element group 159 fork  transition  place  input  bypass 
    -- predecessors 158 
    -- successors 1331 1332 
    -- members (8) 
      -- 	branch_block_stmt_2042/if_stmt_2162_if_link/$exit
      -- 	branch_block_stmt_2042/if_stmt_2162_if_link/if_choice_transition
      -- 	branch_block_stmt_2042/bb_4_bb_7
      -- 	branch_block_stmt_2042/bb_4_bb_7_PhiReq/$entry
      -- 	branch_block_stmt_2042/bb_4_bb_7_PhiReq/phi_stmt_2190/$entry
      -- 	branch_block_stmt_2042/bb_4_bb_7_PhiReq/phi_stmt_2190/phi_stmt_2190_sources/$entry
      -- 	branch_block_stmt_2042/bb_4_bb_7_PhiReq/phi_stmt_2190/phi_stmt_2190_sources/type_cast_2193/$entry
      -- 	branch_block_stmt_2042/bb_4_bb_7_PhiReq/phi_stmt_2190/phi_stmt_2190_sources/type_cast_2193/SplitProtocol/$entry
      -- 
    if_choice_transition_10923_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2162_branch_ack_1, ack => cp_elements(159)); -- 
    -- CP-element group 160 transition  bypass 
    -- predecessors 157 
    -- successors 161 
    -- members (1) 
      -- 	branch_block_stmt_2042/if_stmt_2162_else_link/$entry
      -- 
    cp_elements(160) <= cp_elements(157);
    -- CP-element group 161 transition  place  input  bypass 
    -- predecessors 160 
    -- successors 5 
    -- members (9) 
      -- 	branch_block_stmt_2042/if_stmt_2162_else_link/$exit
      -- 	branch_block_stmt_2042/if_stmt_2162_else_link/else_choice_transition
      -- 	branch_block_stmt_2042/bb_4_bb_5
      -- 	branch_block_stmt_2042/merge_stmt_2168_PhiReqMerge
      -- 	branch_block_stmt_2042/bb_4_bb_5_PhiReq/$entry
      -- 	branch_block_stmt_2042/bb_4_bb_5_PhiReq/$exit
      -- 	branch_block_stmt_2042/merge_stmt_2168_PhiAck/$entry
      -- 	branch_block_stmt_2042/merge_stmt_2168_PhiAck/$exit
      -- 	branch_block_stmt_2042/merge_stmt_2168_PhiAck/dummy
      -- 
    else_choice_transition_10927_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2162_branch_ack_0, ack => cp_elements(161)); -- 
    -- CP-element group 162 fork  transition  bypass 
    -- predecessors 5 
    -- successors 163 164 
    -- members (1) 
      -- 	branch_block_stmt_2042/assign_stmt_2174/$entry
      -- 
    cp_elements(162) <= cp_elements(5);
    -- CP-element group 163 transition  output  bypass 
    -- predecessors 162 
    -- successors 166 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_2174/SGT_f32_u1_2173_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_2174/SGT_f32_u1_2173_Update/$entry
      -- 	branch_block_stmt_2042/assign_stmt_2174/SGT_f32_u1_2173_Update/cr
      -- 
    cp_elements(163) <= cp_elements(162);
    cr_10949_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(163), ack => SGT_f32_u1_2173_inst_req_1); -- 
    -- CP-element group 164 transition  output  bypass 
    -- predecessors 162 
    -- successors 165 
    -- members (7) 
      -- 	branch_block_stmt_2042/assign_stmt_2174/SGT_f32_u1_2173_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_2174/R_iNsTr_17_2170_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_2174/R_iNsTr_17_2170_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2174/R_iNsTr_17_2170_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_2174/R_iNsTr_17_2170_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2174/SGT_f32_u1_2173_Sample/$entry
      -- 	branch_block_stmt_2042/assign_stmt_2174/SGT_f32_u1_2173_Sample/rr
      -- 
    cp_elements(164) <= cp_elements(162);
    rr_10944_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(164), ack => SGT_f32_u1_2173_inst_req_0); -- 
    -- CP-element group 165 transition  input  bypass 
    -- predecessors 164 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_2174/SGT_f32_u1_2173_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2174/SGT_f32_u1_2173_Sample/$exit
      -- 	branch_block_stmt_2042/assign_stmt_2174/SGT_f32_u1_2173_Sample/ra
      -- 
    ra_10945_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => SGT_f32_u1_2173_inst_ack_0, ack => cp_elements(165)); -- 
    -- CP-element group 166 branch  transition  place  input  bypass 
    -- predecessors 163 
    -- successors 167 168 
    -- members (6) 
      -- 	branch_block_stmt_2042/assign_stmt_2174__exit__
      -- 	branch_block_stmt_2042/if_stmt_2175__entry__
      -- 	branch_block_stmt_2042/assign_stmt_2174/$exit
      -- 	branch_block_stmt_2042/assign_stmt_2174/SGT_f32_u1_2173_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2174/SGT_f32_u1_2173_Update/$exit
      -- 	branch_block_stmt_2042/assign_stmt_2174/SGT_f32_u1_2173_Update/ca
      -- 
    ca_10950_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => SGT_f32_u1_2173_inst_ack_1, ack => cp_elements(166)); -- 
    -- CP-element group 167 transition  place  dead  bypass 
    -- predecessors 166 
    -- successors 6 
    -- members (8) 
      -- 	branch_block_stmt_2042/if_stmt_2175__exit__
      -- 	branch_block_stmt_2042/merge_stmt_2181__entry__
      -- 	branch_block_stmt_2042/if_stmt_2175_dead_link/$entry
      -- 	branch_block_stmt_2042/if_stmt_2175_dead_link/$exit
      -- 	branch_block_stmt_2042/if_stmt_2175_dead_link/dead_transition
      -- 	branch_block_stmt_2042/merge_stmt_2181_dead_link/$entry
      -- 	branch_block_stmt_2042/merge_stmt_2181_dead_link/$exit
      -- 	branch_block_stmt_2042/merge_stmt_2181_dead_link/dead_transition
      -- 
    cp_elements(167) <= false;
    -- CP-element group 168 transition  output  bypass 
    -- predecessors 166 
    -- successors 169 
    -- members (3) 
      -- 	branch_block_stmt_2042/if_stmt_2175_eval_test/$entry
      -- 	branch_block_stmt_2042/if_stmt_2175_eval_test/$exit
      -- 	branch_block_stmt_2042/if_stmt_2175_eval_test/branch_req
      -- 
    cp_elements(168) <= cp_elements(166);
    branch_req_10958_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(168), ack => if_stmt_2175_branch_req_0); -- 
    -- CP-element group 169 branch  place  bypass 
    -- predecessors 168 
    -- successors 170 172 
    -- members (1) 
      -- 	branch_block_stmt_2042/R_iNsTr_25_2176_place
      -- 
    cp_elements(169) <= cp_elements(168);
    -- CP-element group 170 transition  bypass 
    -- predecessors 169 
    -- successors 171 
    -- members (1) 
      -- 	branch_block_stmt_2042/if_stmt_2175_if_link/$entry
      -- 
    cp_elements(170) <= cp_elements(169);
    -- CP-element group 171 fork  transition  place  input  bypass 
    -- predecessors 170 
    -- successors 1334 1335 
    -- members (8) 
      -- 	branch_block_stmt_2042/if_stmt_2175_if_link/$exit
      -- 	branch_block_stmt_2042/if_stmt_2175_if_link/if_choice_transition
      -- 	branch_block_stmt_2042/bb_5_bb_7
      -- 	branch_block_stmt_2042/bb_5_bb_7_PhiReq/$entry
      -- 	branch_block_stmt_2042/bb_5_bb_7_PhiReq/phi_stmt_2190/$entry
      -- 	branch_block_stmt_2042/bb_5_bb_7_PhiReq/phi_stmt_2190/phi_stmt_2190_sources/$entry
      -- 	branch_block_stmt_2042/bb_5_bb_7_PhiReq/phi_stmt_2190/phi_stmt_2190_sources/type_cast_2193/$entry
      -- 	branch_block_stmt_2042/bb_5_bb_7_PhiReq/phi_stmt_2190/phi_stmt_2190_sources/type_cast_2193/SplitProtocol/$entry
      -- 
    if_choice_transition_10963_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2175_branch_ack_1, ack => cp_elements(171)); -- 
    -- CP-element group 172 transition  bypass 
    -- predecessors 169 
    -- successors 173 
    -- members (1) 
      -- 	branch_block_stmt_2042/if_stmt_2175_else_link/$entry
      -- 
    cp_elements(172) <= cp_elements(169);
    -- CP-element group 173 transition  place  input  bypass 
    -- predecessors 172 
    -- successors 6 
    -- members (9) 
      -- 	branch_block_stmt_2042/if_stmt_2175_else_link/$exit
      -- 	branch_block_stmt_2042/if_stmt_2175_else_link/else_choice_transition
      -- 	branch_block_stmt_2042/bb_5_bb_6
      -- 	branch_block_stmt_2042/merge_stmt_2181_PhiReqMerge
      -- 	branch_block_stmt_2042/bb_5_bb_6_PhiReq/$entry
      -- 	branch_block_stmt_2042/bb_5_bb_6_PhiReq/$exit
      -- 	branch_block_stmt_2042/merge_stmt_2181_PhiAck/$entry
      -- 	branch_block_stmt_2042/merge_stmt_2181_PhiAck/$exit
      -- 	branch_block_stmt_2042/merge_stmt_2181_PhiAck/dummy
      -- 
    else_choice_transition_10967_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2175_branch_ack_0, ack => cp_elements(173)); -- 
    -- CP-element group 174 fork  transition  bypass 
    -- predecessors 6 
    -- successors 175 176 
    -- members (1) 
      -- 	branch_block_stmt_2042/assign_stmt_2187/$entry
      -- 
    cp_elements(174) <= cp_elements(6);
    -- CP-element group 175 transition  output  bypass 
    -- predecessors 174 
    -- successors 178 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_2187/MUL_f32_f32_2186_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_2187/MUL_f32_f32_2186_Update/$entry
      -- 	branch_block_stmt_2042/assign_stmt_2187/MUL_f32_f32_2186_Update/cr
      -- 
    cp_elements(175) <= cp_elements(174);
    cr_10989_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(175), ack => MUL_f32_f32_2186_inst_req_1); -- 
    -- CP-element group 176 transition  output  bypass 
    -- predecessors 174 
    -- successors 177 
    -- members (7) 
      -- 	branch_block_stmt_2042/assign_stmt_2187/MUL_f32_f32_2186_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_2187/R_iNsTr_17_2183_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_2187/R_iNsTr_17_2183_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2187/R_iNsTr_17_2183_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_2187/R_iNsTr_17_2183_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2187/MUL_f32_f32_2186_Sample/$entry
      -- 	branch_block_stmt_2042/assign_stmt_2187/MUL_f32_f32_2186_Sample/rr
      -- 
    cp_elements(176) <= cp_elements(174);
    rr_10984_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(176), ack => MUL_f32_f32_2186_inst_req_0); -- 
    -- CP-element group 177 transition  input  bypass 
    -- predecessors 176 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_2187/MUL_f32_f32_2186_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2187/MUL_f32_f32_2186_Sample/$exit
      -- 	branch_block_stmt_2042/assign_stmt_2187/MUL_f32_f32_2186_Sample/ra
      -- 
    ra_10985_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => MUL_f32_f32_2186_inst_ack_0, ack => cp_elements(177)); -- 
    -- CP-element group 178 fork  transition  place  input  bypass 
    -- predecessors 175 
    -- successors 1337 1339 
    -- members (11) 
      -- 	branch_block_stmt_2042/assign_stmt_2187__exit__
      -- 	branch_block_stmt_2042/bb_6_bb_7
      -- 	branch_block_stmt_2042/assign_stmt_2187/$exit
      -- 	branch_block_stmt_2042/assign_stmt_2187/MUL_f32_f32_2186_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2187/MUL_f32_f32_2186_Update/$exit
      -- 	branch_block_stmt_2042/assign_stmt_2187/MUL_f32_f32_2186_Update/ca
      -- 	branch_block_stmt_2042/bb_6_bb_7_PhiReq/$entry
      -- 	branch_block_stmt_2042/bb_6_bb_7_PhiReq/phi_stmt_2190/$entry
      -- 	branch_block_stmt_2042/bb_6_bb_7_PhiReq/phi_stmt_2190/phi_stmt_2190_sources/$entry
      -- 	branch_block_stmt_2042/bb_6_bb_7_PhiReq/phi_stmt_2190/phi_stmt_2190_sources/type_cast_2193/$entry
      -- 	branch_block_stmt_2042/bb_6_bb_7_PhiReq/phi_stmt_2190/phi_stmt_2190_sources/type_cast_2193/SplitProtocol/$entry
      -- 
    ca_10990_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => MUL_f32_f32_2186_inst_ack_1, ack => cp_elements(178)); -- 
    -- CP-element group 179 fork  transition  bypass 
    -- predecessors 1344 
    -- successors 180 181 184 
    -- members (1) 
      -- 	branch_block_stmt_2042/assign_stmt_2204_to_assign_stmt_2210/$entry
      -- 
    cp_elements(179) <= cp_elements(1344);
    -- CP-element group 180 transition  output  bypass 
    -- predecessors 179 
    -- successors 183 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_2204_to_assign_stmt_2210/type_cast_2203_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_2204_to_assign_stmt_2210/type_cast_2203_Update/$entry
      -- 	branch_block_stmt_2042/assign_stmt_2204_to_assign_stmt_2210/type_cast_2203_Update/cr
      -- 
    cp_elements(180) <= cp_elements(179);
    cr_11010_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(180), ack => type_cast_2203_inst_req_1); -- 
    -- CP-element group 181 transition  output  bypass 
    -- predecessors 179 
    -- successors 182 
    -- members (7) 
      -- 	branch_block_stmt_2042/assign_stmt_2204_to_assign_stmt_2210/type_cast_2203_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_2204_to_assign_stmt_2210/R_iNsTr_8_2202_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_2204_to_assign_stmt_2210/R_iNsTr_8_2202_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2204_to_assign_stmt_2210/R_iNsTr_8_2202_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_2204_to_assign_stmt_2210/R_iNsTr_8_2202_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2204_to_assign_stmt_2210/type_cast_2203_Sample/$entry
      -- 	branch_block_stmt_2042/assign_stmt_2204_to_assign_stmt_2210/type_cast_2203_Sample/rr
      -- 
    cp_elements(181) <= cp_elements(179);
    rr_11005_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(181), ack => type_cast_2203_inst_req_0); -- 
    -- CP-element group 182 transition  input  bypass 
    -- predecessors 181 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_2204_to_assign_stmt_2210/type_cast_2203_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2204_to_assign_stmt_2210/type_cast_2203_Sample/$exit
      -- 	branch_block_stmt_2042/assign_stmt_2204_to_assign_stmt_2210/type_cast_2203_Sample/ra
      -- 
    ra_11006_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2203_inst_ack_0, ack => cp_elements(182)); -- 
    -- CP-element group 183 transition  input  output  bypass 
    -- predecessors 180 
    -- successors 185 
    -- members (10) 
      -- 	branch_block_stmt_2042/assign_stmt_2204_to_assign_stmt_2210/type_cast_2203_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2204_to_assign_stmt_2210/type_cast_2203_Update/$exit
      -- 	branch_block_stmt_2042/assign_stmt_2204_to_assign_stmt_2210/type_cast_2203_Update/ca
      -- 	branch_block_stmt_2042/assign_stmt_2204_to_assign_stmt_2210/SGT_f64_u1_2209_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_2204_to_assign_stmt_2210/R_iNsTr_22_2206_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_2204_to_assign_stmt_2210/R_iNsTr_22_2206_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2204_to_assign_stmt_2210/R_iNsTr_22_2206_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_2204_to_assign_stmt_2210/R_iNsTr_22_2206_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2204_to_assign_stmt_2210/SGT_f64_u1_2209_Sample/$entry
      -- 	branch_block_stmt_2042/assign_stmt_2204_to_assign_stmt_2210/SGT_f64_u1_2209_Sample/rr
      -- 
    ca_11011_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2203_inst_ack_1, ack => cp_elements(183)); -- 
    rr_11023_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(183), ack => SGT_f64_u1_2209_inst_req_0); -- 
    -- CP-element group 184 transition  output  bypass 
    -- predecessors 179 
    -- successors 186 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_2204_to_assign_stmt_2210/SGT_f64_u1_2209_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_2204_to_assign_stmt_2210/SGT_f64_u1_2209_Update/$entry
      -- 	branch_block_stmt_2042/assign_stmt_2204_to_assign_stmt_2210/SGT_f64_u1_2209_Update/cr
      -- 
    cp_elements(184) <= cp_elements(179);
    cr_11028_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(184), ack => SGT_f64_u1_2209_inst_req_1); -- 
    -- CP-element group 185 transition  input  bypass 
    -- predecessors 183 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_2204_to_assign_stmt_2210/SGT_f64_u1_2209_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2204_to_assign_stmt_2210/SGT_f64_u1_2209_Sample/$exit
      -- 	branch_block_stmt_2042/assign_stmt_2204_to_assign_stmt_2210/SGT_f64_u1_2209_Sample/ra
      -- 
    ra_11024_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => SGT_f64_u1_2209_inst_ack_0, ack => cp_elements(185)); -- 
    -- CP-element group 186 branch  transition  place  input  bypass 
    -- predecessors 184 
    -- successors 187 188 
    -- members (6) 
      -- 	branch_block_stmt_2042/assign_stmt_2204_to_assign_stmt_2210__exit__
      -- 	branch_block_stmt_2042/if_stmt_2211__entry__
      -- 	branch_block_stmt_2042/assign_stmt_2204_to_assign_stmt_2210/$exit
      -- 	branch_block_stmt_2042/assign_stmt_2204_to_assign_stmt_2210/SGT_f64_u1_2209_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2204_to_assign_stmt_2210/SGT_f64_u1_2209_Update/$exit
      -- 	branch_block_stmt_2042/assign_stmt_2204_to_assign_stmt_2210/SGT_f64_u1_2209_Update/ca
      -- 
    ca_11029_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => SGT_f64_u1_2209_inst_ack_1, ack => cp_elements(186)); -- 
    -- CP-element group 187 transition  place  dead  bypass 
    -- predecessors 186 
    -- successors 7 
    -- members (8) 
      -- 	branch_block_stmt_2042/if_stmt_2211__exit__
      -- 	branch_block_stmt_2042/merge_stmt_2217__entry__
      -- 	branch_block_stmt_2042/if_stmt_2211_dead_link/$entry
      -- 	branch_block_stmt_2042/if_stmt_2211_dead_link/$exit
      -- 	branch_block_stmt_2042/if_stmt_2211_dead_link/dead_transition
      -- 	branch_block_stmt_2042/merge_stmt_2217_dead_link/$entry
      -- 	branch_block_stmt_2042/merge_stmt_2217_dead_link/$exit
      -- 	branch_block_stmt_2042/merge_stmt_2217_dead_link/dead_transition
      -- 
    cp_elements(187) <= false;
    -- CP-element group 188 transition  output  bypass 
    -- predecessors 186 
    -- successors 189 
    -- members (3) 
      -- 	branch_block_stmt_2042/if_stmt_2211_eval_test/$entry
      -- 	branch_block_stmt_2042/if_stmt_2211_eval_test/$exit
      -- 	branch_block_stmt_2042/if_stmt_2211_eval_test/branch_req
      -- 
    cp_elements(188) <= cp_elements(186);
    branch_req_11037_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(188), ack => if_stmt_2211_branch_req_0); -- 
    -- CP-element group 189 branch  place  bypass 
    -- predecessors 188 
    -- successors 190 192 
    -- members (1) 
      -- 	branch_block_stmt_2042/R_iNsTr_23_2212_place
      -- 
    cp_elements(189) <= cp_elements(188);
    -- CP-element group 190 transition  bypass 
    -- predecessors 189 
    -- successors 191 
    -- members (1) 
      -- 	branch_block_stmt_2042/if_stmt_2211_if_link/$entry
      -- 
    cp_elements(190) <= cp_elements(189);
    -- CP-element group 191 transition  place  input  bypass 
    -- predecessors 190 
    -- successors 7 
    -- members (9) 
      -- 	branch_block_stmt_2042/if_stmt_2211_if_link/$exit
      -- 	branch_block_stmt_2042/if_stmt_2211_if_link/if_choice_transition
      -- 	branch_block_stmt_2042/bb_7_bb_8
      -- 	branch_block_stmt_2042/merge_stmt_2217_PhiReqMerge
      -- 	branch_block_stmt_2042/bb_7_bb_8_PhiReq/$entry
      -- 	branch_block_stmt_2042/bb_7_bb_8_PhiReq/$exit
      -- 	branch_block_stmt_2042/merge_stmt_2217_PhiAck/$entry
      -- 	branch_block_stmt_2042/merge_stmt_2217_PhiAck/$exit
      -- 	branch_block_stmt_2042/merge_stmt_2217_PhiAck/dummy
      -- 
    if_choice_transition_11042_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2211_branch_ack_1, ack => cp_elements(191)); -- 
    -- CP-element group 192 transition  bypass 
    -- predecessors 189 
    -- successors 193 
    -- members (1) 
      -- 	branch_block_stmt_2042/if_stmt_2211_else_link/$entry
      -- 
    cp_elements(192) <= cp_elements(189);
    -- CP-element group 193 fork  transition  place  input  bypass 
    -- predecessors 192 
    -- successors 1375 1379 1383 
    -- members (6) 
      -- 	branch_block_stmt_2042/if_stmt_2211_else_link/$exit
      -- 	branch_block_stmt_2042/if_stmt_2211_else_link/else_choice_transition
      -- 	branch_block_stmt_2042/bb_7_bb_13
      -- 	branch_block_stmt_2042/bb_7_bb_13_PhiReq/$entry
      -- 	branch_block_stmt_2042/bb_7_bb_13_PhiReq/phi_stmt_2304/$entry
      -- 	branch_block_stmt_2042/bb_7_bb_13_PhiReq/phi_stmt_2304/phi_stmt_2304_sources/$entry
      -- 
    else_choice_transition_11046_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2211_branch_ack_0, ack => cp_elements(193)); -- 
    -- CP-element group 194 fork  transition  bypass 
    -- predecessors 7 
    -- successors 195 196 
    -- members (1) 
      -- 	branch_block_stmt_2042/assign_stmt_2223/$entry
      -- 
    cp_elements(194) <= cp_elements(7);
    -- CP-element group 195 transition  output  bypass 
    -- predecessors 194 
    -- successors 198 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_2223/SGT_f64_u1_2222_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_2223/SGT_f64_u1_2222_Update/$entry
      -- 	branch_block_stmt_2042/assign_stmt_2223/SGT_f64_u1_2222_Update/cr
      -- 
    cp_elements(195) <= cp_elements(194);
    cr_11068_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(195), ack => SGT_f64_u1_2222_inst_req_1); -- 
    -- CP-element group 196 transition  output  bypass 
    -- predecessors 194 
    -- successors 197 
    -- members (7) 
      -- 	branch_block_stmt_2042/assign_stmt_2223/SGT_f64_u1_2222_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_2223/R_iNsTr_22_2219_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_2223/R_iNsTr_22_2219_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2223/R_iNsTr_22_2219_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_2223/R_iNsTr_22_2219_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2223/SGT_f64_u1_2222_Sample/$entry
      -- 	branch_block_stmt_2042/assign_stmt_2223/SGT_f64_u1_2222_Sample/rr
      -- 
    cp_elements(196) <= cp_elements(194);
    rr_11063_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(196), ack => SGT_f64_u1_2222_inst_req_0); -- 
    -- CP-element group 197 transition  input  bypass 
    -- predecessors 196 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_2223/SGT_f64_u1_2222_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2223/SGT_f64_u1_2222_Sample/$exit
      -- 	branch_block_stmt_2042/assign_stmt_2223/SGT_f64_u1_2222_Sample/ra
      -- 
    ra_11064_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => SGT_f64_u1_2222_inst_ack_0, ack => cp_elements(197)); -- 
    -- CP-element group 198 branch  transition  place  input  bypass 
    -- predecessors 195 
    -- successors 199 200 
    -- members (6) 
      -- 	branch_block_stmt_2042/assign_stmt_2223__exit__
      -- 	branch_block_stmt_2042/if_stmt_2224__entry__
      -- 	branch_block_stmt_2042/assign_stmt_2223/$exit
      -- 	branch_block_stmt_2042/assign_stmt_2223/SGT_f64_u1_2222_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2223/SGT_f64_u1_2222_Update/$exit
      -- 	branch_block_stmt_2042/assign_stmt_2223/SGT_f64_u1_2222_Update/ca
      -- 
    ca_11069_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => SGT_f64_u1_2222_inst_ack_1, ack => cp_elements(198)); -- 
    -- CP-element group 199 transition  place  dead  bypass 
    -- predecessors 198 
    -- successors 8 
    -- members (8) 
      -- 	branch_block_stmt_2042/if_stmt_2224__exit__
      -- 	branch_block_stmt_2042/merge_stmt_2230__entry__
      -- 	branch_block_stmt_2042/if_stmt_2224_dead_link/$entry
      -- 	branch_block_stmt_2042/if_stmt_2224_dead_link/$exit
      -- 	branch_block_stmt_2042/if_stmt_2224_dead_link/dead_transition
      -- 	branch_block_stmt_2042/merge_stmt_2230_dead_link/$entry
      -- 	branch_block_stmt_2042/merge_stmt_2230_dead_link/$exit
      -- 	branch_block_stmt_2042/merge_stmt_2230_dead_link/dead_transition
      -- 
    cp_elements(199) <= false;
    -- CP-element group 200 transition  output  bypass 
    -- predecessors 198 
    -- successors 201 
    -- members (3) 
      -- 	branch_block_stmt_2042/if_stmt_2224_eval_test/$entry
      -- 	branch_block_stmt_2042/if_stmt_2224_eval_test/$exit
      -- 	branch_block_stmt_2042/if_stmt_2224_eval_test/branch_req
      -- 
    cp_elements(200) <= cp_elements(198);
    branch_req_11077_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(200), ack => if_stmt_2224_branch_req_0); -- 
    -- CP-element group 201 branch  place  bypass 
    -- predecessors 200 
    -- successors 202 204 
    -- members (1) 
      -- 	branch_block_stmt_2042/R_iNsTr_28_2225_place
      -- 
    cp_elements(201) <= cp_elements(200);
    -- CP-element group 202 transition  bypass 
    -- predecessors 201 
    -- successors 203 
    -- members (1) 
      -- 	branch_block_stmt_2042/if_stmt_2224_if_link/$entry
      -- 
    cp_elements(202) <= cp_elements(201);
    -- CP-element group 203 transition  place  input  bypass 
    -- predecessors 202 
    -- successors 217 
    -- members (11) 
      -- 	branch_block_stmt_2042/merge_stmt_2250__exit__
      -- 	branch_block_stmt_2042/assign_stmt_2256__entry__
      -- 	branch_block_stmt_2042/if_stmt_2224_if_link/$exit
      -- 	branch_block_stmt_2042/if_stmt_2224_if_link/if_choice_transition
      -- 	branch_block_stmt_2042/bb_8_bb_10
      -- 	branch_block_stmt_2042/merge_stmt_2250_PhiReqMerge
      -- 	branch_block_stmt_2042/bb_8_bb_10_PhiReq/$entry
      -- 	branch_block_stmt_2042/bb_8_bb_10_PhiReq/$exit
      -- 	branch_block_stmt_2042/merge_stmt_2250_PhiAck/$entry
      -- 	branch_block_stmt_2042/merge_stmt_2250_PhiAck/$exit
      -- 	branch_block_stmt_2042/merge_stmt_2250_PhiAck/dummy
      -- 
    if_choice_transition_11082_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2224_branch_ack_1, ack => cp_elements(203)); -- 
    -- CP-element group 204 transition  bypass 
    -- predecessors 201 
    -- successors 205 
    -- members (1) 
      -- 	branch_block_stmt_2042/if_stmt_2224_else_link/$entry
      -- 
    cp_elements(204) <= cp_elements(201);
    -- CP-element group 205 transition  place  input  bypass 
    -- predecessors 204 
    -- successors 8 
    -- members (9) 
      -- 	branch_block_stmt_2042/if_stmt_2224_else_link/$exit
      -- 	branch_block_stmt_2042/if_stmt_2224_else_link/else_choice_transition
      -- 	branch_block_stmt_2042/bb_8_bb_9
      -- 	branch_block_stmt_2042/merge_stmt_2230_PhiReqMerge
      -- 	branch_block_stmt_2042/bb_8_bb_9_PhiReq/$entry
      -- 	branch_block_stmt_2042/bb_8_bb_9_PhiReq/$exit
      -- 	branch_block_stmt_2042/merge_stmt_2230_PhiAck/$entry
      -- 	branch_block_stmt_2042/merge_stmt_2230_PhiAck/$exit
      -- 	branch_block_stmt_2042/merge_stmt_2230_PhiAck/dummy
      -- 
    else_choice_transition_11086_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2224_branch_ack_0, ack => cp_elements(205)); -- 
    -- CP-element group 206 fork  transition  bypass 
    -- predecessors 8 
    -- successors 207 208 211 214 
    -- members (1) 
      -- 	branch_block_stmt_2042/assign_stmt_2236_to_assign_stmt_2248/$entry
      -- 
    cp_elements(206) <= cp_elements(8);
    -- CP-element group 207 transition  output  bypass 
    -- predecessors 206 
    -- successors 210 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_2236_to_assign_stmt_2248/MUL_f32_f32_2235_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_2236_to_assign_stmt_2248/MUL_f32_f32_2235_Update/$entry
      -- 	branch_block_stmt_2042/assign_stmt_2236_to_assign_stmt_2248/MUL_f32_f32_2235_Update/cr
      -- 
    cp_elements(207) <= cp_elements(206);
    cr_11108_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(207), ack => MUL_f32_f32_2235_inst_req_1); -- 
    -- CP-element group 208 transition  output  bypass 
    -- predecessors 206 
    -- successors 209 
    -- members (7) 
      -- 	branch_block_stmt_2042/assign_stmt_2236_to_assign_stmt_2248/MUL_f32_f32_2235_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_2236_to_assign_stmt_2248/R_iNsTr_8_2232_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_2236_to_assign_stmt_2248/R_iNsTr_8_2232_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2236_to_assign_stmt_2248/R_iNsTr_8_2232_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_2236_to_assign_stmt_2248/R_iNsTr_8_2232_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2236_to_assign_stmt_2248/MUL_f32_f32_2235_Sample/$entry
      -- 	branch_block_stmt_2042/assign_stmt_2236_to_assign_stmt_2248/MUL_f32_f32_2235_Sample/rr
      -- 
    cp_elements(208) <= cp_elements(206);
    rr_11103_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(208), ack => MUL_f32_f32_2235_inst_req_0); -- 
    -- CP-element group 209 transition  input  bypass 
    -- predecessors 208 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_2236_to_assign_stmt_2248/MUL_f32_f32_2235_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2236_to_assign_stmt_2248/MUL_f32_f32_2235_Sample/$exit
      -- 	branch_block_stmt_2042/assign_stmt_2236_to_assign_stmt_2248/MUL_f32_f32_2235_Sample/ra
      -- 
    ra_11104_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => MUL_f32_f32_2235_inst_ack_0, ack => cp_elements(209)); -- 
    -- CP-element group 210 transition  input  output  bypass 
    -- predecessors 207 
    -- successors 212 
    -- members (10) 
      -- 	branch_block_stmt_2042/assign_stmt_2236_to_assign_stmt_2248/MUL_f32_f32_2235_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2236_to_assign_stmt_2248/MUL_f32_f32_2235_Update/$exit
      -- 	branch_block_stmt_2042/assign_stmt_2236_to_assign_stmt_2248/MUL_f32_f32_2235_Update/ca
      -- 	branch_block_stmt_2042/assign_stmt_2236_to_assign_stmt_2248/ADD_f32_f32_2241_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_2236_to_assign_stmt_2248/R_iNsTr_38_2238_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_2236_to_assign_stmt_2248/R_iNsTr_38_2238_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2236_to_assign_stmt_2248/R_iNsTr_38_2238_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_2236_to_assign_stmt_2248/R_iNsTr_38_2238_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2236_to_assign_stmt_2248/ADD_f32_f32_2241_Sample/$entry
      -- 	branch_block_stmt_2042/assign_stmt_2236_to_assign_stmt_2248/ADD_f32_f32_2241_Sample/rr
      -- 
    ca_11109_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => MUL_f32_f32_2235_inst_ack_1, ack => cp_elements(210)); -- 
    rr_11121_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(210), ack => ADD_f32_f32_2241_inst_req_0); -- 
    -- CP-element group 211 transition  output  bypass 
    -- predecessors 206 
    -- successors 213 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_2236_to_assign_stmt_2248/ADD_f32_f32_2241_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_2236_to_assign_stmt_2248/ADD_f32_f32_2241_Update/$entry
      -- 	branch_block_stmt_2042/assign_stmt_2236_to_assign_stmt_2248/ADD_f32_f32_2241_Update/cr
      -- 
    cp_elements(211) <= cp_elements(206);
    cr_11126_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(211), ack => ADD_f32_f32_2241_inst_req_1); -- 
    -- CP-element group 212 transition  input  bypass 
    -- predecessors 210 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_2236_to_assign_stmt_2248/ADD_f32_f32_2241_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2236_to_assign_stmt_2248/ADD_f32_f32_2241_Sample/$exit
      -- 	branch_block_stmt_2042/assign_stmt_2236_to_assign_stmt_2248/ADD_f32_f32_2241_Sample/ra
      -- 
    ra_11122_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_f32_f32_2241_inst_ack_0, ack => cp_elements(212)); -- 
    -- CP-element group 213 transition  input  output  bypass 
    -- predecessors 211 
    -- successors 215 
    -- members (10) 
      -- 	branch_block_stmt_2042/assign_stmt_2236_to_assign_stmt_2248/ADD_f32_f32_2241_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2236_to_assign_stmt_2248/ADD_f32_f32_2241_Update/$exit
      -- 	branch_block_stmt_2042/assign_stmt_2236_to_assign_stmt_2248/ADD_f32_f32_2241_Update/ca
      -- 	branch_block_stmt_2042/assign_stmt_2236_to_assign_stmt_2248/MUL_f32_f32_2247_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_2236_to_assign_stmt_2248/R_iNsTr_39_2244_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_2236_to_assign_stmt_2248/R_iNsTr_39_2244_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2236_to_assign_stmt_2248/R_iNsTr_39_2244_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_2236_to_assign_stmt_2248/R_iNsTr_39_2244_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2236_to_assign_stmt_2248/MUL_f32_f32_2247_Sample/$entry
      -- 	branch_block_stmt_2042/assign_stmt_2236_to_assign_stmt_2248/MUL_f32_f32_2247_Sample/rr
      -- 
    ca_11127_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_f32_f32_2241_inst_ack_1, ack => cp_elements(213)); -- 
    rr_11139_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(213), ack => MUL_f32_f32_2247_inst_req_0); -- 
    -- CP-element group 214 transition  output  bypass 
    -- predecessors 206 
    -- successors 216 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_2236_to_assign_stmt_2248/MUL_f32_f32_2247_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_2236_to_assign_stmt_2248/MUL_f32_f32_2247_Update/$entry
      -- 	branch_block_stmt_2042/assign_stmt_2236_to_assign_stmt_2248/MUL_f32_f32_2247_Update/cr
      -- 
    cp_elements(214) <= cp_elements(206);
    cr_11144_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(214), ack => MUL_f32_f32_2247_inst_req_1); -- 
    -- CP-element group 215 transition  input  bypass 
    -- predecessors 213 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_2236_to_assign_stmt_2248/MUL_f32_f32_2247_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2236_to_assign_stmt_2248/MUL_f32_f32_2247_Sample/$exit
      -- 	branch_block_stmt_2042/assign_stmt_2236_to_assign_stmt_2248/MUL_f32_f32_2247_Sample/ra
      -- 
    ra_11140_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => MUL_f32_f32_2247_inst_ack_0, ack => cp_elements(215)); -- 
    -- CP-element group 216 fork  transition  place  input  bypass 
    -- predecessors 214 
    -- successors 1388 1394 1398 
    -- members (9) 
      -- 	branch_block_stmt_2042/assign_stmt_2236_to_assign_stmt_2248__exit__
      -- 	branch_block_stmt_2042/bb_9_bb_13
      -- 	branch_block_stmt_2042/assign_stmt_2236_to_assign_stmt_2248/$exit
      -- 	branch_block_stmt_2042/assign_stmt_2236_to_assign_stmt_2248/MUL_f32_f32_2247_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2236_to_assign_stmt_2248/MUL_f32_f32_2247_Update/$exit
      -- 	branch_block_stmt_2042/assign_stmt_2236_to_assign_stmt_2248/MUL_f32_f32_2247_Update/ca
      -- 	branch_block_stmt_2042/bb_9_bb_13_PhiReq/$entry
      -- 	branch_block_stmt_2042/bb_9_bb_13_PhiReq/phi_stmt_2304/$entry
      -- 	branch_block_stmt_2042/bb_9_bb_13_PhiReq/phi_stmt_2304/phi_stmt_2304_sources/$entry
      -- 
    ca_11145_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => MUL_f32_f32_2247_inst_ack_1, ack => cp_elements(216)); -- 
    -- CP-element group 217 fork  transition  bypass 
    -- predecessors 203 
    -- successors 218 219 
    -- members (1) 
      -- 	branch_block_stmt_2042/assign_stmt_2256/$entry
      -- 
    cp_elements(217) <= cp_elements(203);
    -- CP-element group 218 transition  output  bypass 
    -- predecessors 217 
    -- successors 221 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_2256/SGT_f64_u1_2255_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_2256/SGT_f64_u1_2255_Update/$entry
      -- 	branch_block_stmt_2042/assign_stmt_2256/SGT_f64_u1_2255_Update/cr
      -- 
    cp_elements(218) <= cp_elements(217);
    cr_11165_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(218), ack => SGT_f64_u1_2255_inst_req_1); -- 
    -- CP-element group 219 transition  output  bypass 
    -- predecessors 217 
    -- successors 220 
    -- members (7) 
      -- 	branch_block_stmt_2042/assign_stmt_2256/SGT_f64_u1_2255_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_2256/R_iNsTr_22_2252_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_2256/R_iNsTr_22_2252_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2256/R_iNsTr_22_2252_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_2256/R_iNsTr_22_2252_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2256/SGT_f64_u1_2255_Sample/$entry
      -- 	branch_block_stmt_2042/assign_stmt_2256/SGT_f64_u1_2255_Sample/rr
      -- 
    cp_elements(219) <= cp_elements(217);
    rr_11160_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(219), ack => SGT_f64_u1_2255_inst_req_0); -- 
    -- CP-element group 220 transition  input  bypass 
    -- predecessors 219 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_2256/SGT_f64_u1_2255_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2256/SGT_f64_u1_2255_Sample/$exit
      -- 	branch_block_stmt_2042/assign_stmt_2256/SGT_f64_u1_2255_Sample/ra
      -- 
    ra_11161_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => SGT_f64_u1_2255_inst_ack_0, ack => cp_elements(220)); -- 
    -- CP-element group 221 branch  transition  place  input  bypass 
    -- predecessors 218 
    -- successors 222 223 
    -- members (6) 
      -- 	branch_block_stmt_2042/assign_stmt_2256__exit__
      -- 	branch_block_stmt_2042/if_stmt_2257__entry__
      -- 	branch_block_stmt_2042/assign_stmt_2256/$exit
      -- 	branch_block_stmt_2042/assign_stmt_2256/SGT_f64_u1_2255_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2256/SGT_f64_u1_2255_Update/$exit
      -- 	branch_block_stmt_2042/assign_stmt_2256/SGT_f64_u1_2255_Update/ca
      -- 
    ca_11166_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => SGT_f64_u1_2255_inst_ack_1, ack => cp_elements(221)); -- 
    -- CP-element group 222 transition  place  dead  bypass 
    -- predecessors 221 
    -- successors 9 
    -- members (8) 
      -- 	branch_block_stmt_2042/if_stmt_2257__exit__
      -- 	branch_block_stmt_2042/merge_stmt_2263__entry__
      -- 	branch_block_stmt_2042/if_stmt_2257_dead_link/$entry
      -- 	branch_block_stmt_2042/if_stmt_2257_dead_link/$exit
      -- 	branch_block_stmt_2042/if_stmt_2257_dead_link/dead_transition
      -- 	branch_block_stmt_2042/merge_stmt_2263_dead_link/$entry
      -- 	branch_block_stmt_2042/merge_stmt_2263_dead_link/$exit
      -- 	branch_block_stmt_2042/merge_stmt_2263_dead_link/dead_transition
      -- 
    cp_elements(222) <= false;
    -- CP-element group 223 transition  output  bypass 
    -- predecessors 221 
    -- successors 224 
    -- members (3) 
      -- 	branch_block_stmt_2042/if_stmt_2257_eval_test/$entry
      -- 	branch_block_stmt_2042/if_stmt_2257_eval_test/$exit
      -- 	branch_block_stmt_2042/if_stmt_2257_eval_test/branch_req
      -- 
    cp_elements(223) <= cp_elements(221);
    branch_req_11174_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(223), ack => if_stmt_2257_branch_req_0); -- 
    -- CP-element group 224 branch  place  bypass 
    -- predecessors 223 
    -- successors 225 227 
    -- members (1) 
      -- 	branch_block_stmt_2042/R_iNsTr_36_2258_place
      -- 
    cp_elements(224) <= cp_elements(223);
    -- CP-element group 225 transition  bypass 
    -- predecessors 224 
    -- successors 226 
    -- members (1) 
      -- 	branch_block_stmt_2042/if_stmt_2257_if_link/$entry
      -- 
    cp_elements(225) <= cp_elements(224);
    -- CP-element group 226 transition  place  input  bypass 
    -- predecessors 225 
    -- successors 240 
    -- members (11) 
      -- 	branch_block_stmt_2042/merge_stmt_2283__exit__
      -- 	branch_block_stmt_2042/assign_stmt_2289_to_assign_stmt_2301__entry__
      -- 	branch_block_stmt_2042/if_stmt_2257_if_link/$exit
      -- 	branch_block_stmt_2042/if_stmt_2257_if_link/if_choice_transition
      -- 	branch_block_stmt_2042/bb_10_bb_12
      -- 	branch_block_stmt_2042/merge_stmt_2283_PhiReqMerge
      -- 	branch_block_stmt_2042/bb_10_bb_12_PhiReq/$entry
      -- 	branch_block_stmt_2042/bb_10_bb_12_PhiReq/$exit
      -- 	branch_block_stmt_2042/merge_stmt_2283_PhiAck/$entry
      -- 	branch_block_stmt_2042/merge_stmt_2283_PhiAck/$exit
      -- 	branch_block_stmt_2042/merge_stmt_2283_PhiAck/dummy
      -- 
    if_choice_transition_11179_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2257_branch_ack_1, ack => cp_elements(226)); -- 
    -- CP-element group 227 transition  bypass 
    -- predecessors 224 
    -- successors 228 
    -- members (1) 
      -- 	branch_block_stmt_2042/if_stmt_2257_else_link/$entry
      -- 
    cp_elements(227) <= cp_elements(224);
    -- CP-element group 228 transition  place  input  bypass 
    -- predecessors 227 
    -- successors 9 
    -- members (9) 
      -- 	branch_block_stmt_2042/if_stmt_2257_else_link/$exit
      -- 	branch_block_stmt_2042/if_stmt_2257_else_link/else_choice_transition
      -- 	branch_block_stmt_2042/bb_10_bb_11
      -- 	branch_block_stmt_2042/merge_stmt_2263_PhiReqMerge
      -- 	branch_block_stmt_2042/bb_10_bb_11_PhiReq/$entry
      -- 	branch_block_stmt_2042/bb_10_bb_11_PhiReq/$exit
      -- 	branch_block_stmt_2042/merge_stmt_2263_PhiAck/$entry
      -- 	branch_block_stmt_2042/merge_stmt_2263_PhiAck/$exit
      -- 	branch_block_stmt_2042/merge_stmt_2263_PhiAck/dummy
      -- 
    else_choice_transition_11183_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2257_branch_ack_0, ack => cp_elements(228)); -- 
    -- CP-element group 229 fork  transition  bypass 
    -- predecessors 9 
    -- successors 230 231 234 237 
    -- members (1) 
      -- 	branch_block_stmt_2042/assign_stmt_2269_to_assign_stmt_2281/$entry
      -- 
    cp_elements(229) <= cp_elements(9);
    -- CP-element group 230 transition  output  bypass 
    -- predecessors 229 
    -- successors 233 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_2269_to_assign_stmt_2281/MUL_f32_f32_2268_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_2269_to_assign_stmt_2281/MUL_f32_f32_2268_Update/$entry
      -- 	branch_block_stmt_2042/assign_stmt_2269_to_assign_stmt_2281/MUL_f32_f32_2268_Update/cr
      -- 
    cp_elements(230) <= cp_elements(229);
    cr_11205_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(230), ack => MUL_f32_f32_2268_inst_req_1); -- 
    -- CP-element group 231 transition  output  bypass 
    -- predecessors 229 
    -- successors 232 
    -- members (7) 
      -- 	branch_block_stmt_2042/assign_stmt_2269_to_assign_stmt_2281/MUL_f32_f32_2268_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_2269_to_assign_stmt_2281/R_iNsTr_8_2265_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_2269_to_assign_stmt_2281/R_iNsTr_8_2265_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2269_to_assign_stmt_2281/R_iNsTr_8_2265_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_2269_to_assign_stmt_2281/R_iNsTr_8_2265_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2269_to_assign_stmt_2281/MUL_f32_f32_2268_Sample/$entry
      -- 	branch_block_stmt_2042/assign_stmt_2269_to_assign_stmt_2281/MUL_f32_f32_2268_Sample/rr
      -- 
    cp_elements(231) <= cp_elements(229);
    rr_11200_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(231), ack => MUL_f32_f32_2268_inst_req_0); -- 
    -- CP-element group 232 transition  input  bypass 
    -- predecessors 231 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_2269_to_assign_stmt_2281/MUL_f32_f32_2268_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2269_to_assign_stmt_2281/MUL_f32_f32_2268_Sample/$exit
      -- 	branch_block_stmt_2042/assign_stmt_2269_to_assign_stmt_2281/MUL_f32_f32_2268_Sample/ra
      -- 
    ra_11201_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => MUL_f32_f32_2268_inst_ack_0, ack => cp_elements(232)); -- 
    -- CP-element group 233 transition  input  output  bypass 
    -- predecessors 230 
    -- successors 235 
    -- members (10) 
      -- 	branch_block_stmt_2042/assign_stmt_2269_to_assign_stmt_2281/MUL_f32_f32_2268_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2269_to_assign_stmt_2281/MUL_f32_f32_2268_Update/$exit
      -- 	branch_block_stmt_2042/assign_stmt_2269_to_assign_stmt_2281/MUL_f32_f32_2268_Update/ca
      -- 	branch_block_stmt_2042/assign_stmt_2269_to_assign_stmt_2281/ADD_f32_f32_2274_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_2269_to_assign_stmt_2281/R_iNsTr_55_2271_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_2269_to_assign_stmt_2281/R_iNsTr_55_2271_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2269_to_assign_stmt_2281/R_iNsTr_55_2271_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_2269_to_assign_stmt_2281/R_iNsTr_55_2271_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2269_to_assign_stmt_2281/ADD_f32_f32_2274_Sample/$entry
      -- 	branch_block_stmt_2042/assign_stmt_2269_to_assign_stmt_2281/ADD_f32_f32_2274_Sample/rr
      -- 
    ca_11206_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => MUL_f32_f32_2268_inst_ack_1, ack => cp_elements(233)); -- 
    rr_11218_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(233), ack => ADD_f32_f32_2274_inst_req_0); -- 
    -- CP-element group 234 transition  output  bypass 
    -- predecessors 229 
    -- successors 236 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_2269_to_assign_stmt_2281/ADD_f32_f32_2274_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_2269_to_assign_stmt_2281/ADD_f32_f32_2274_Update/$entry
      -- 	branch_block_stmt_2042/assign_stmt_2269_to_assign_stmt_2281/ADD_f32_f32_2274_Update/cr
      -- 
    cp_elements(234) <= cp_elements(229);
    cr_11223_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(234), ack => ADD_f32_f32_2274_inst_req_1); -- 
    -- CP-element group 235 transition  input  bypass 
    -- predecessors 233 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_2269_to_assign_stmt_2281/ADD_f32_f32_2274_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2269_to_assign_stmt_2281/ADD_f32_f32_2274_Sample/$exit
      -- 	branch_block_stmt_2042/assign_stmt_2269_to_assign_stmt_2281/ADD_f32_f32_2274_Sample/ra
      -- 
    ra_11219_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_f32_f32_2274_inst_ack_0, ack => cp_elements(235)); -- 
    -- CP-element group 236 transition  input  output  bypass 
    -- predecessors 234 
    -- successors 238 
    -- members (10) 
      -- 	branch_block_stmt_2042/assign_stmt_2269_to_assign_stmt_2281/ADD_f32_f32_2274_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2269_to_assign_stmt_2281/ADD_f32_f32_2274_Update/$exit
      -- 	branch_block_stmt_2042/assign_stmt_2269_to_assign_stmt_2281/ADD_f32_f32_2274_Update/ca
      -- 	branch_block_stmt_2042/assign_stmt_2269_to_assign_stmt_2281/MUL_f32_f32_2280_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_2269_to_assign_stmt_2281/R_iNsTr_56_2277_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_2269_to_assign_stmt_2281/R_iNsTr_56_2277_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2269_to_assign_stmt_2281/R_iNsTr_56_2277_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_2269_to_assign_stmt_2281/R_iNsTr_56_2277_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2269_to_assign_stmt_2281/MUL_f32_f32_2280_Sample/$entry
      -- 	branch_block_stmt_2042/assign_stmt_2269_to_assign_stmt_2281/MUL_f32_f32_2280_Sample/rr
      -- 
    ca_11224_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_f32_f32_2274_inst_ack_1, ack => cp_elements(236)); -- 
    rr_11236_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(236), ack => MUL_f32_f32_2280_inst_req_0); -- 
    -- CP-element group 237 transition  output  bypass 
    -- predecessors 229 
    -- successors 239 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_2269_to_assign_stmt_2281/MUL_f32_f32_2280_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_2269_to_assign_stmt_2281/MUL_f32_f32_2280_Update/$entry
      -- 	branch_block_stmt_2042/assign_stmt_2269_to_assign_stmt_2281/MUL_f32_f32_2280_Update/cr
      -- 
    cp_elements(237) <= cp_elements(229);
    cr_11241_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(237), ack => MUL_f32_f32_2280_inst_req_1); -- 
    -- CP-element group 238 transition  input  bypass 
    -- predecessors 236 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_2269_to_assign_stmt_2281/MUL_f32_f32_2280_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2269_to_assign_stmt_2281/MUL_f32_f32_2280_Sample/$exit
      -- 	branch_block_stmt_2042/assign_stmt_2269_to_assign_stmt_2281/MUL_f32_f32_2280_Sample/ra
      -- 
    ra_11237_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => MUL_f32_f32_2280_inst_ack_0, ack => cp_elements(238)); -- 
    -- CP-element group 239 fork  transition  place  input  bypass 
    -- predecessors 237 
    -- successors 1345 1349 1355 
    -- members (9) 
      -- 	branch_block_stmt_2042/assign_stmt_2269_to_assign_stmt_2281__exit__
      -- 	branch_block_stmt_2042/bb_11_bb_13
      -- 	branch_block_stmt_2042/assign_stmt_2269_to_assign_stmt_2281/$exit
      -- 	branch_block_stmt_2042/assign_stmt_2269_to_assign_stmt_2281/MUL_f32_f32_2280_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2269_to_assign_stmt_2281/MUL_f32_f32_2280_Update/$exit
      -- 	branch_block_stmt_2042/assign_stmt_2269_to_assign_stmt_2281/MUL_f32_f32_2280_Update/ca
      -- 	branch_block_stmt_2042/bb_11_bb_13_PhiReq/$entry
      -- 	branch_block_stmt_2042/bb_11_bb_13_PhiReq/phi_stmt_2304/$entry
      -- 	branch_block_stmt_2042/bb_11_bb_13_PhiReq/phi_stmt_2304/phi_stmt_2304_sources/$entry
      -- 
    ca_11242_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => MUL_f32_f32_2280_inst_ack_1, ack => cp_elements(239)); -- 
    -- CP-element group 240 fork  transition  bypass 
    -- predecessors 226 
    -- successors 241 242 245 248 
    -- members (1) 
      -- 	branch_block_stmt_2042/assign_stmt_2289_to_assign_stmt_2301/$entry
      -- 
    cp_elements(240) <= cp_elements(226);
    -- CP-element group 241 transition  output  bypass 
    -- predecessors 240 
    -- successors 244 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_2289_to_assign_stmt_2301/MUL_f32_f32_2288_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_2289_to_assign_stmt_2301/MUL_f32_f32_2288_Update/$entry
      -- 	branch_block_stmt_2042/assign_stmt_2289_to_assign_stmt_2301/MUL_f32_f32_2288_Update/cr
      -- 
    cp_elements(241) <= cp_elements(240);
    cr_11262_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(241), ack => MUL_f32_f32_2288_inst_req_1); -- 
    -- CP-element group 242 transition  output  bypass 
    -- predecessors 240 
    -- successors 243 
    -- members (7) 
      -- 	branch_block_stmt_2042/assign_stmt_2289_to_assign_stmt_2301/MUL_f32_f32_2288_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_2289_to_assign_stmt_2301/R_iNsTr_8_2285_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_2289_to_assign_stmt_2301/R_iNsTr_8_2285_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2289_to_assign_stmt_2301/R_iNsTr_8_2285_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_2289_to_assign_stmt_2301/R_iNsTr_8_2285_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2289_to_assign_stmt_2301/MUL_f32_f32_2288_Sample/$entry
      -- 	branch_block_stmt_2042/assign_stmt_2289_to_assign_stmt_2301/MUL_f32_f32_2288_Sample/rr
      -- 
    cp_elements(242) <= cp_elements(240);
    rr_11257_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(242), ack => MUL_f32_f32_2288_inst_req_0); -- 
    -- CP-element group 243 transition  input  bypass 
    -- predecessors 242 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_2289_to_assign_stmt_2301/MUL_f32_f32_2288_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2289_to_assign_stmt_2301/MUL_f32_f32_2288_Sample/$exit
      -- 	branch_block_stmt_2042/assign_stmt_2289_to_assign_stmt_2301/MUL_f32_f32_2288_Sample/ra
      -- 
    ra_11258_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => MUL_f32_f32_2288_inst_ack_0, ack => cp_elements(243)); -- 
    -- CP-element group 244 transition  input  output  bypass 
    -- predecessors 241 
    -- successors 246 
    -- members (10) 
      -- 	branch_block_stmt_2042/assign_stmt_2289_to_assign_stmt_2301/MUL_f32_f32_2288_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2289_to_assign_stmt_2301/MUL_f32_f32_2288_Update/$exit
      -- 	branch_block_stmt_2042/assign_stmt_2289_to_assign_stmt_2301/MUL_f32_f32_2288_Update/ca
      -- 	branch_block_stmt_2042/assign_stmt_2289_to_assign_stmt_2301/ADD_f32_f32_2294_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_2289_to_assign_stmt_2301/R_iNsTr_51_2291_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_2289_to_assign_stmt_2301/R_iNsTr_51_2291_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2289_to_assign_stmt_2301/R_iNsTr_51_2291_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_2289_to_assign_stmt_2301/R_iNsTr_51_2291_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2289_to_assign_stmt_2301/ADD_f32_f32_2294_Sample/$entry
      -- 	branch_block_stmt_2042/assign_stmt_2289_to_assign_stmt_2301/ADD_f32_f32_2294_Sample/rr
      -- 
    ca_11263_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => MUL_f32_f32_2288_inst_ack_1, ack => cp_elements(244)); -- 
    rr_11275_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(244), ack => ADD_f32_f32_2294_inst_req_0); -- 
    -- CP-element group 245 transition  output  bypass 
    -- predecessors 240 
    -- successors 247 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_2289_to_assign_stmt_2301/ADD_f32_f32_2294_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_2289_to_assign_stmt_2301/ADD_f32_f32_2294_Update/$entry
      -- 	branch_block_stmt_2042/assign_stmt_2289_to_assign_stmt_2301/ADD_f32_f32_2294_Update/cr
      -- 
    cp_elements(245) <= cp_elements(240);
    cr_11280_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(245), ack => ADD_f32_f32_2294_inst_req_1); -- 
    -- CP-element group 246 transition  input  bypass 
    -- predecessors 244 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_2289_to_assign_stmt_2301/ADD_f32_f32_2294_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2289_to_assign_stmt_2301/ADD_f32_f32_2294_Sample/$exit
      -- 	branch_block_stmt_2042/assign_stmt_2289_to_assign_stmt_2301/ADD_f32_f32_2294_Sample/ra
      -- 
    ra_11276_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_f32_f32_2294_inst_ack_0, ack => cp_elements(246)); -- 
    -- CP-element group 247 transition  input  output  bypass 
    -- predecessors 245 
    -- successors 249 
    -- members (10) 
      -- 	branch_block_stmt_2042/assign_stmt_2289_to_assign_stmt_2301/ADD_f32_f32_2294_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2289_to_assign_stmt_2301/ADD_f32_f32_2294_Update/$exit
      -- 	branch_block_stmt_2042/assign_stmt_2289_to_assign_stmt_2301/ADD_f32_f32_2294_Update/ca
      -- 	branch_block_stmt_2042/assign_stmt_2289_to_assign_stmt_2301/MUL_f32_f32_2300_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_2289_to_assign_stmt_2301/R_iNsTr_52_2297_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_2289_to_assign_stmt_2301/R_iNsTr_52_2297_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2289_to_assign_stmt_2301/R_iNsTr_52_2297_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_2289_to_assign_stmt_2301/R_iNsTr_52_2297_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2289_to_assign_stmt_2301/MUL_f32_f32_2300_Sample/$entry
      -- 	branch_block_stmt_2042/assign_stmt_2289_to_assign_stmt_2301/MUL_f32_f32_2300_Sample/rr
      -- 
    ca_11281_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_f32_f32_2294_inst_ack_1, ack => cp_elements(247)); -- 
    rr_11293_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(247), ack => MUL_f32_f32_2300_inst_req_0); -- 
    -- CP-element group 248 transition  output  bypass 
    -- predecessors 240 
    -- successors 250 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_2289_to_assign_stmt_2301/MUL_f32_f32_2300_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_2289_to_assign_stmt_2301/MUL_f32_f32_2300_Update/$entry
      -- 	branch_block_stmt_2042/assign_stmt_2289_to_assign_stmt_2301/MUL_f32_f32_2300_Update/cr
      -- 
    cp_elements(248) <= cp_elements(240);
    cr_11298_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(248), ack => MUL_f32_f32_2300_inst_req_1); -- 
    -- CP-element group 249 transition  input  bypass 
    -- predecessors 247 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_2289_to_assign_stmt_2301/MUL_f32_f32_2300_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2289_to_assign_stmt_2301/MUL_f32_f32_2300_Sample/$exit
      -- 	branch_block_stmt_2042/assign_stmt_2289_to_assign_stmt_2301/MUL_f32_f32_2300_Sample/ra
      -- 
    ra_11294_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => MUL_f32_f32_2300_inst_ack_0, ack => cp_elements(249)); -- 
    -- CP-element group 250 fork  transition  place  input  bypass 
    -- predecessors 248 
    -- successors 1360 1364 1368 
    -- members (9) 
      -- 	branch_block_stmt_2042/assign_stmt_2289_to_assign_stmt_2301__exit__
      -- 	branch_block_stmt_2042/bb_12_bb_13
      -- 	branch_block_stmt_2042/assign_stmt_2289_to_assign_stmt_2301/$exit
      -- 	branch_block_stmt_2042/assign_stmt_2289_to_assign_stmt_2301/MUL_f32_f32_2300_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2289_to_assign_stmt_2301/MUL_f32_f32_2300_Update/$exit
      -- 	branch_block_stmt_2042/assign_stmt_2289_to_assign_stmt_2301/MUL_f32_f32_2300_Update/ca
      -- 	branch_block_stmt_2042/bb_12_bb_13_PhiReq/$entry
      -- 	branch_block_stmt_2042/bb_12_bb_13_PhiReq/phi_stmt_2304/$entry
      -- 	branch_block_stmt_2042/bb_12_bb_13_PhiReq/phi_stmt_2304/phi_stmt_2304_sources/$entry
      -- 
    ca_11299_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => MUL_f32_f32_2300_inst_ack_1, ack => cp_elements(250)); -- 
    -- CP-element group 251 fork  transition  bypass 
    -- predecessors 1405 
    -- successors 252 253 256 257 261 264 268 
    -- members (1) 
      -- 	branch_block_stmt_2042/assign_stmt_2321_to_assign_stmt_2342/$entry
      -- 
    cp_elements(251) <= cp_elements(1405);
    -- CP-element group 252 transition  output  bypass 
    -- predecessors 251 
    -- successors 255 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_2321_to_assign_stmt_2342/MUL_f32_f32_2320_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_2321_to_assign_stmt_2342/MUL_f32_f32_2320_Update/$entry
      -- 	branch_block_stmt_2042/assign_stmt_2321_to_assign_stmt_2342/MUL_f32_f32_2320_Update/cr
      -- 
    cp_elements(252) <= cp_elements(251);
    cr_11319_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(252), ack => MUL_f32_f32_2320_inst_req_1); -- 
    -- CP-element group 253 transition  output  bypass 
    -- predecessors 251 
    -- successors 254 
    -- members (7) 
      -- 	branch_block_stmt_2042/assign_stmt_2321_to_assign_stmt_2342/MUL_f32_f32_2320_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_2321_to_assign_stmt_2342/R_iNsTr_2_2317_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_2321_to_assign_stmt_2342/R_iNsTr_2_2317_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2321_to_assign_stmt_2342/R_iNsTr_2_2317_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_2321_to_assign_stmt_2342/R_iNsTr_2_2317_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2321_to_assign_stmt_2342/MUL_f32_f32_2320_Sample/$entry
      -- 	branch_block_stmt_2042/assign_stmt_2321_to_assign_stmt_2342/MUL_f32_f32_2320_Sample/rr
      -- 
    cp_elements(253) <= cp_elements(251);
    rr_11314_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(253), ack => MUL_f32_f32_2320_inst_req_0); -- 
    -- CP-element group 254 transition  input  bypass 
    -- predecessors 253 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_2321_to_assign_stmt_2342/MUL_f32_f32_2320_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2321_to_assign_stmt_2342/MUL_f32_f32_2320_Sample/$exit
      -- 	branch_block_stmt_2042/assign_stmt_2321_to_assign_stmt_2342/MUL_f32_f32_2320_Sample/ra
      -- 
    ra_11315_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => MUL_f32_f32_2320_inst_ack_0, ack => cp_elements(254)); -- 
    -- CP-element group 255 transition  input  bypass 
    -- predecessors 252 
    -- successors 260 
    -- members (7) 
      -- 	branch_block_stmt_2042/assign_stmt_2321_to_assign_stmt_2342/MUL_f32_f32_2320_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2321_to_assign_stmt_2342/MUL_f32_f32_2320_Update/$exit
      -- 	branch_block_stmt_2042/assign_stmt_2321_to_assign_stmt_2342/MUL_f32_f32_2320_Update/ca
      -- 	branch_block_stmt_2042/assign_stmt_2321_to_assign_stmt_2342/R_iNsTr_30_2330_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_2321_to_assign_stmt_2342/R_iNsTr_30_2330_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2321_to_assign_stmt_2342/R_iNsTr_30_2330_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_2321_to_assign_stmt_2342/R_iNsTr_30_2330_update_completed_
      -- 
    ca_11320_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => MUL_f32_f32_2320_inst_ack_1, ack => cp_elements(255)); -- 
    -- CP-element group 256 transition  output  bypass 
    -- predecessors 251 
    -- successors 259 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_2321_to_assign_stmt_2342/MUL_f32_f32_2326_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_2321_to_assign_stmt_2342/MUL_f32_f32_2326_Update/$entry
      -- 	branch_block_stmt_2042/assign_stmt_2321_to_assign_stmt_2342/MUL_f32_f32_2326_Update/cr
      -- 
    cp_elements(256) <= cp_elements(251);
    cr_11337_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(256), ack => MUL_f32_f32_2326_inst_req_1); -- 
    -- CP-element group 257 transition  output  bypass 
    -- predecessors 251 
    -- successors 258 
    -- members (7) 
      -- 	branch_block_stmt_2042/assign_stmt_2321_to_assign_stmt_2342/MUL_f32_f32_2326_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_2321_to_assign_stmt_2342/R_flux_rotor_prevx_x0_2323_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_2321_to_assign_stmt_2342/R_flux_rotor_prevx_x0_2323_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2321_to_assign_stmt_2342/R_flux_rotor_prevx_x0_2323_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_2321_to_assign_stmt_2342/R_flux_rotor_prevx_x0_2323_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2321_to_assign_stmt_2342/MUL_f32_f32_2326_Sample/$entry
      -- 	branch_block_stmt_2042/assign_stmt_2321_to_assign_stmt_2342/MUL_f32_f32_2326_Sample/rr
      -- 
    cp_elements(257) <= cp_elements(251);
    rr_11332_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(257), ack => MUL_f32_f32_2326_inst_req_0); -- 
    -- CP-element group 258 transition  input  bypass 
    -- predecessors 257 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_2321_to_assign_stmt_2342/MUL_f32_f32_2326_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2321_to_assign_stmt_2342/MUL_f32_f32_2326_Sample/$exit
      -- 	branch_block_stmt_2042/assign_stmt_2321_to_assign_stmt_2342/MUL_f32_f32_2326_Sample/ra
      -- 
    ra_11333_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => MUL_f32_f32_2326_inst_ack_0, ack => cp_elements(258)); -- 
    -- CP-element group 259 transition  input  bypass 
    -- predecessors 256 
    -- successors 260 
    -- members (7) 
      -- 	branch_block_stmt_2042/assign_stmt_2321_to_assign_stmt_2342/MUL_f32_f32_2326_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2321_to_assign_stmt_2342/MUL_f32_f32_2326_Update/$exit
      -- 	branch_block_stmt_2042/assign_stmt_2321_to_assign_stmt_2342/MUL_f32_f32_2326_Update/ca
      -- 	branch_block_stmt_2042/assign_stmt_2321_to_assign_stmt_2342/R_iNsTr_31_2329_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_2321_to_assign_stmt_2342/R_iNsTr_31_2329_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2321_to_assign_stmt_2342/R_iNsTr_31_2329_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_2321_to_assign_stmt_2342/R_iNsTr_31_2329_update_completed_
      -- 
    ca_11338_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => MUL_f32_f32_2326_inst_ack_1, ack => cp_elements(259)); -- 
    -- CP-element group 260 join  transition  output  bypass 
    -- predecessors 255 259 
    -- successors 262 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_2321_to_assign_stmt_2342/ADD_f32_f32_2331_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_2321_to_assign_stmt_2342/ADD_f32_f32_2331_Sample/$entry
      -- 	branch_block_stmt_2042/assign_stmt_2321_to_assign_stmt_2342/ADD_f32_f32_2331_Sample/rr
      -- 
    cp_element_group_260: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 20) := "cp_element_group_260"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(255) & cp_elements(259);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(260), clk => clk, reset => reset); --
    end block;
    rr_11354_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(260), ack => ADD_f32_f32_2331_inst_req_0); -- 
    -- CP-element group 261 transition  output  bypass 
    -- predecessors 251 
    -- successors 263 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_2321_to_assign_stmt_2342/ADD_f32_f32_2331_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_2321_to_assign_stmt_2342/ADD_f32_f32_2331_Update/$entry
      -- 	branch_block_stmt_2042/assign_stmt_2321_to_assign_stmt_2342/ADD_f32_f32_2331_Update/cr
      -- 
    cp_elements(261) <= cp_elements(251);
    cr_11359_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(261), ack => ADD_f32_f32_2331_inst_req_1); -- 
    -- CP-element group 262 transition  input  bypass 
    -- predecessors 260 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_2321_to_assign_stmt_2342/ADD_f32_f32_2331_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2321_to_assign_stmt_2342/ADD_f32_f32_2331_Sample/$exit
      -- 	branch_block_stmt_2042/assign_stmt_2321_to_assign_stmt_2342/ADD_f32_f32_2331_Sample/ra
      -- 
    ra_11355_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_f32_f32_2331_inst_ack_0, ack => cp_elements(262)); -- 
    -- CP-element group 263 fork  transition  input  bypass 
    -- predecessors 261 
    -- successors 265 269 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_2321_to_assign_stmt_2342/ADD_f32_f32_2331_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2321_to_assign_stmt_2342/ADD_f32_f32_2331_Update/$exit
      -- 	branch_block_stmt_2042/assign_stmt_2321_to_assign_stmt_2342/ADD_f32_f32_2331_Update/ca
      -- 
    ca_11360_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_f32_f32_2331_inst_ack_1, ack => cp_elements(263)); -- 
    -- CP-element group 264 transition  output  bypass 
    -- predecessors 251 
    -- successors 267 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_2321_to_assign_stmt_2342/type_cast_2335_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_2321_to_assign_stmt_2342/type_cast_2335_Update/$entry
      -- 	branch_block_stmt_2042/assign_stmt_2321_to_assign_stmt_2342/type_cast_2335_Update/cr
      -- 
    cp_elements(264) <= cp_elements(251);
    cr_11377_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(264), ack => type_cast_2335_inst_req_1); -- 
    -- CP-element group 265 transition  output  bypass 
    -- predecessors 263 
    -- successors 266 
    -- members (7) 
      -- 	branch_block_stmt_2042/assign_stmt_2321_to_assign_stmt_2342/type_cast_2335_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_2321_to_assign_stmt_2342/R_iNsTr_32_2334_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_2321_to_assign_stmt_2342/R_iNsTr_32_2334_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2321_to_assign_stmt_2342/R_iNsTr_32_2334_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_2321_to_assign_stmt_2342/R_iNsTr_32_2334_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2321_to_assign_stmt_2342/type_cast_2335_Sample/$entry
      -- 	branch_block_stmt_2042/assign_stmt_2321_to_assign_stmt_2342/type_cast_2335_Sample/rr
      -- 
    cp_elements(265) <= cp_elements(263);
    rr_11372_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(265), ack => type_cast_2335_inst_req_0); -- 
    -- CP-element group 266 transition  input  bypass 
    -- predecessors 265 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_2321_to_assign_stmt_2342/type_cast_2335_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2321_to_assign_stmt_2342/type_cast_2335_Sample/$exit
      -- 	branch_block_stmt_2042/assign_stmt_2321_to_assign_stmt_2342/type_cast_2335_Sample/ra
      -- 
    ra_11373_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2335_inst_ack_0, ack => cp_elements(266)); -- 
    -- CP-element group 267 transition  input  bypass 
    -- predecessors 264 
    -- successors 272 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_2321_to_assign_stmt_2342/type_cast_2335_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2321_to_assign_stmt_2342/type_cast_2335_Update/$exit
      -- 	branch_block_stmt_2042/assign_stmt_2321_to_assign_stmt_2342/type_cast_2335_Update/ca
      -- 
    ca_11378_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2335_inst_ack_1, ack => cp_elements(267)); -- 
    -- CP-element group 268 transition  output  bypass 
    -- predecessors 251 
    -- successors 271 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_2321_to_assign_stmt_2342/EQ_f32_u1_2341_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_2321_to_assign_stmt_2342/EQ_f32_u1_2341_Update/$entry
      -- 	branch_block_stmt_2042/assign_stmt_2321_to_assign_stmt_2342/EQ_f32_u1_2341_Update/cr
      -- 
    cp_elements(268) <= cp_elements(251);
    cr_11395_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(268), ack => EQ_f32_u1_2341_inst_req_1); -- 
    -- CP-element group 269 transition  output  bypass 
    -- predecessors 263 
    -- successors 270 
    -- members (7) 
      -- 	branch_block_stmt_2042/assign_stmt_2321_to_assign_stmt_2342/EQ_f32_u1_2341_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_2321_to_assign_stmt_2342/R_iNsTr_32_2338_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_2321_to_assign_stmt_2342/R_iNsTr_32_2338_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2321_to_assign_stmt_2342/R_iNsTr_32_2338_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_2321_to_assign_stmt_2342/R_iNsTr_32_2338_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2321_to_assign_stmt_2342/EQ_f32_u1_2341_Sample/$entry
      -- 	branch_block_stmt_2042/assign_stmt_2321_to_assign_stmt_2342/EQ_f32_u1_2341_Sample/rr
      -- 
    cp_elements(269) <= cp_elements(263);
    rr_11390_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(269), ack => EQ_f32_u1_2341_inst_req_0); -- 
    -- CP-element group 270 transition  input  bypass 
    -- predecessors 269 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_2321_to_assign_stmt_2342/EQ_f32_u1_2341_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2321_to_assign_stmt_2342/EQ_f32_u1_2341_Sample/$exit
      -- 	branch_block_stmt_2042/assign_stmt_2321_to_assign_stmt_2342/EQ_f32_u1_2341_Sample/ra
      -- 
    ra_11391_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_f32_u1_2341_inst_ack_0, ack => cp_elements(270)); -- 
    -- CP-element group 271 transition  input  bypass 
    -- predecessors 268 
    -- successors 272 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_2321_to_assign_stmt_2342/EQ_f32_u1_2341_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2321_to_assign_stmt_2342/EQ_f32_u1_2341_Update/$exit
      -- 	branch_block_stmt_2042/assign_stmt_2321_to_assign_stmt_2342/EQ_f32_u1_2341_Update/ca
      -- 
    ca_11396_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_f32_u1_2341_inst_ack_1, ack => cp_elements(271)); -- 
    -- CP-element group 272 join  transition  bypass 
    -- predecessors 267 271 
    -- successors 10 
    -- members (1) 
      -- 	branch_block_stmt_2042/assign_stmt_2321_to_assign_stmt_2342/$exit
      -- 
    cp_element_group_272: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 20) := "cp_element_group_272"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(267) & cp_elements(271);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(272), clk => clk, reset => reset); --
    end block;
    -- CP-element group 273 transition  place  dead  bypass 
    -- predecessors 10 
    -- successors 11 
    -- members (8) 
      -- 	branch_block_stmt_2042/if_stmt_2343__exit__
      -- 	branch_block_stmt_2042/merge_stmt_2349__entry__
      -- 	branch_block_stmt_2042/if_stmt_2343_dead_link/$entry
      -- 	branch_block_stmt_2042/if_stmt_2343_dead_link/$exit
      -- 	branch_block_stmt_2042/if_stmt_2343_dead_link/dead_transition
      -- 	branch_block_stmt_2042/merge_stmt_2349_dead_link/$entry
      -- 	branch_block_stmt_2042/merge_stmt_2349_dead_link/$exit
      -- 	branch_block_stmt_2042/merge_stmt_2349_dead_link/dead_transition
      -- 
    cp_elements(273) <= false;
    -- CP-element group 274 transition  output  bypass 
    -- predecessors 10 
    -- successors 275 
    -- members (3) 
      -- 	branch_block_stmt_2042/if_stmt_2343_eval_test/$entry
      -- 	branch_block_stmt_2042/if_stmt_2343_eval_test/$exit
      -- 	branch_block_stmt_2042/if_stmt_2343_eval_test/branch_req
      -- 
    cp_elements(274) <= cp_elements(10);
    branch_req_11404_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(274), ack => if_stmt_2343_branch_req_0); -- 
    -- CP-element group 275 branch  place  bypass 
    -- predecessors 274 
    -- successors 276 278 
    -- members (1) 
      -- 	branch_block_stmt_2042/R_iNsTr_33_2344_place
      -- 
    cp_elements(275) <= cp_elements(274);
    -- CP-element group 276 transition  bypass 
    -- predecessors 275 
    -- successors 277 
    -- members (1) 
      -- 	branch_block_stmt_2042/if_stmt_2343_if_link/$entry
      -- 
    cp_elements(276) <= cp_elements(275);
    -- CP-element group 277 fork  transition  place  input  bypass 
    -- predecessors 276 
    -- successors 1651 1652 
    -- members (8) 
      -- 	branch_block_stmt_2042/if_stmt_2343_if_link/if_choice_transition
      -- 	branch_block_stmt_2042/if_stmt_2343_if_link/$exit
      -- 	branch_block_stmt_2042/bb_13_rotor_flux_calcx_xexit
      -- 	branch_block_stmt_2042/bb_13_rotor_flux_calcx_xexit_PhiReq/$entry
      -- 	branch_block_stmt_2042/bb_13_rotor_flux_calcx_xexit_PhiReq/phi_stmt_2683/$entry
      -- 	branch_block_stmt_2042/bb_13_rotor_flux_calcx_xexit_PhiReq/phi_stmt_2683/phi_stmt_2683_sources/$entry
      -- 	branch_block_stmt_2042/bb_13_rotor_flux_calcx_xexit_PhiReq/phi_stmt_2683/phi_stmt_2683_sources/type_cast_2686/$entry
      -- 	branch_block_stmt_2042/bb_13_rotor_flux_calcx_xexit_PhiReq/phi_stmt_2683/phi_stmt_2683_sources/type_cast_2686/SplitProtocol/$entry
      -- 
    if_choice_transition_11409_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2343_branch_ack_1, ack => cp_elements(277)); -- 
    -- CP-element group 278 transition  bypass 
    -- predecessors 275 
    -- successors 279 
    -- members (1) 
      -- 	branch_block_stmt_2042/if_stmt_2343_else_link/$entry
      -- 
    cp_elements(278) <= cp_elements(275);
    -- CP-element group 279 transition  place  input  bypass 
    -- predecessors 278 
    -- successors 11 
    -- members (9) 
      -- 	branch_block_stmt_2042/if_stmt_2343_else_link/else_choice_transition
      -- 	branch_block_stmt_2042/if_stmt_2343_else_link/$exit
      -- 	branch_block_stmt_2042/bb_13_bb_14
      -- 	branch_block_stmt_2042/merge_stmt_2349_PhiReqMerge
      -- 	branch_block_stmt_2042/bb_13_bb_14_PhiReq/$entry
      -- 	branch_block_stmt_2042/bb_13_bb_14_PhiReq/$exit
      -- 	branch_block_stmt_2042/merge_stmt_2349_PhiAck/$entry
      -- 	branch_block_stmt_2042/merge_stmt_2349_PhiAck/$exit
      -- 	branch_block_stmt_2042/merge_stmt_2349_PhiAck/dummy
      -- 
    else_choice_transition_11413_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2343_branch_ack_0, ack => cp_elements(279)); -- 
    -- CP-element group 280 fork  transition  bypass 
    -- predecessors 11 
    -- successors 281 282 285 288 
    -- members (1) 
      -- 	branch_block_stmt_2042/assign_stmt_2355_to_assign_stmt_2367/$entry
      -- 
    cp_elements(280) <= cp_elements(11);
    -- CP-element group 281 transition  output  bypass 
    -- predecessors 280 
    -- successors 284 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_2355_to_assign_stmt_2367/SHL_u32_u32_2354_Update/$entry
      -- 	branch_block_stmt_2042/assign_stmt_2355_to_assign_stmt_2367/SHL_u32_u32_2354_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_2355_to_assign_stmt_2367/SHL_u32_u32_2354_Update/cr
      -- 
    cp_elements(281) <= cp_elements(280);
    cr_11435_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(281), ack => SHL_u32_u32_2354_inst_req_1); -- 
    -- CP-element group 282 transition  output  bypass 
    -- predecessors 280 
    -- successors 283 
    -- members (7) 
      -- 	branch_block_stmt_2042/assign_stmt_2355_to_assign_stmt_2367/SHL_u32_u32_2354_Sample/rr
      -- 	branch_block_stmt_2042/assign_stmt_2355_to_assign_stmt_2367/SHL_u32_u32_2354_Sample/$entry
      -- 	branch_block_stmt_2042/assign_stmt_2355_to_assign_stmt_2367/R_tmp10x_xix_xi30_2351_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2355_to_assign_stmt_2367/R_tmp10x_xix_xi30_2351_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_2355_to_assign_stmt_2367/R_tmp10x_xix_xi30_2351_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2355_to_assign_stmt_2367/R_tmp10x_xix_xi30_2351_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_2355_to_assign_stmt_2367/SHL_u32_u32_2354_sample_start_
      -- 
    cp_elements(282) <= cp_elements(280);
    rr_11430_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(282), ack => SHL_u32_u32_2354_inst_req_0); -- 
    -- CP-element group 283 transition  input  bypass 
    -- predecessors 282 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_2355_to_assign_stmt_2367/SHL_u32_u32_2354_Sample/ra
      -- 	branch_block_stmt_2042/assign_stmt_2355_to_assign_stmt_2367/SHL_u32_u32_2354_Sample/$exit
      -- 	branch_block_stmt_2042/assign_stmt_2355_to_assign_stmt_2367/SHL_u32_u32_2354_sample_completed_
      -- 
    ra_11431_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => SHL_u32_u32_2354_inst_ack_0, ack => cp_elements(283)); -- 
    -- CP-element group 284 transition  input  output  bypass 
    -- predecessors 281 
    -- successors 286 
    -- members (10) 
      -- 	branch_block_stmt_2042/assign_stmt_2355_to_assign_stmt_2367/SHL_u32_u32_2354_Update/ca
      -- 	branch_block_stmt_2042/assign_stmt_2355_to_assign_stmt_2367/AND_u32_u32_2360_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_2355_to_assign_stmt_2367/SHL_u32_u32_2354_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2355_to_assign_stmt_2367/SHL_u32_u32_2354_Update/$exit
      -- 	branch_block_stmt_2042/assign_stmt_2355_to_assign_stmt_2367/AND_u32_u32_2360_Sample/rr
      -- 	branch_block_stmt_2042/assign_stmt_2355_to_assign_stmt_2367/AND_u32_u32_2360_Sample/$entry
      -- 	branch_block_stmt_2042/assign_stmt_2355_to_assign_stmt_2367/R_iNsTr_47_2357_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2355_to_assign_stmt_2367/R_iNsTr_47_2357_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_2355_to_assign_stmt_2367/R_iNsTr_47_2357_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2355_to_assign_stmt_2367/R_iNsTr_47_2357_sample_start_
      -- 
    ca_11436_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => SHL_u32_u32_2354_inst_ack_1, ack => cp_elements(284)); -- 
    rr_11448_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(284), ack => AND_u32_u32_2360_inst_req_0); -- 
    -- CP-element group 285 transition  output  bypass 
    -- predecessors 280 
    -- successors 287 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_2355_to_assign_stmt_2367/AND_u32_u32_2360_Update/cr
      -- 	branch_block_stmt_2042/assign_stmt_2355_to_assign_stmt_2367/AND_u32_u32_2360_Update/$entry
      -- 	branch_block_stmt_2042/assign_stmt_2355_to_assign_stmt_2367/AND_u32_u32_2360_update_start_
      -- 
    cp_elements(285) <= cp_elements(280);
    cr_11453_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(285), ack => AND_u32_u32_2360_inst_req_1); -- 
    -- CP-element group 286 transition  input  bypass 
    -- predecessors 284 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_2355_to_assign_stmt_2367/AND_u32_u32_2360_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2355_to_assign_stmt_2367/AND_u32_u32_2360_Sample/ra
      -- 	branch_block_stmt_2042/assign_stmt_2355_to_assign_stmt_2367/AND_u32_u32_2360_Sample/$exit
      -- 
    ra_11449_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => AND_u32_u32_2360_inst_ack_0, ack => cp_elements(286)); -- 
    -- CP-element group 287 transition  input  output  bypass 
    -- predecessors 285 
    -- successors 289 
    -- members (10) 
      -- 	branch_block_stmt_2042/assign_stmt_2355_to_assign_stmt_2367/OR_u32_u32_2366_Sample/rr
      -- 	branch_block_stmt_2042/assign_stmt_2355_to_assign_stmt_2367/OR_u32_u32_2366_Sample/$entry
      -- 	branch_block_stmt_2042/assign_stmt_2355_to_assign_stmt_2367/R_iNsTr_48_2363_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2355_to_assign_stmt_2367/R_iNsTr_48_2363_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_2355_to_assign_stmt_2367/R_iNsTr_48_2363_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2355_to_assign_stmt_2367/R_iNsTr_48_2363_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_2355_to_assign_stmt_2367/OR_u32_u32_2366_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_2355_to_assign_stmt_2367/AND_u32_u32_2360_Update/ca
      -- 	branch_block_stmt_2042/assign_stmt_2355_to_assign_stmt_2367/AND_u32_u32_2360_Update/$exit
      -- 	branch_block_stmt_2042/assign_stmt_2355_to_assign_stmt_2367/AND_u32_u32_2360_update_completed_
      -- 
    ca_11454_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => AND_u32_u32_2360_inst_ack_1, ack => cp_elements(287)); -- 
    rr_11466_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(287), ack => OR_u32_u32_2366_inst_req_0); -- 
    -- CP-element group 288 transition  output  bypass 
    -- predecessors 280 
    -- successors 290 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_2355_to_assign_stmt_2367/OR_u32_u32_2366_Update/cr
      -- 	branch_block_stmt_2042/assign_stmt_2355_to_assign_stmt_2367/OR_u32_u32_2366_Update/$entry
      -- 	branch_block_stmt_2042/assign_stmt_2355_to_assign_stmt_2367/OR_u32_u32_2366_update_start_
      -- 
    cp_elements(288) <= cp_elements(280);
    cr_11471_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(288), ack => OR_u32_u32_2366_inst_req_1); -- 
    -- CP-element group 289 transition  input  bypass 
    -- predecessors 287 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_2355_to_assign_stmt_2367/OR_u32_u32_2366_Sample/ra
      -- 	branch_block_stmt_2042/assign_stmt_2355_to_assign_stmt_2367/OR_u32_u32_2366_Sample/$exit
      -- 	branch_block_stmt_2042/assign_stmt_2355_to_assign_stmt_2367/OR_u32_u32_2366_sample_completed_
      -- 
    ra_11467_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => OR_u32_u32_2366_inst_ack_0, ack => cp_elements(289)); -- 
    -- CP-element group 290 transition  place  input  bypass 
    -- predecessors 288 
    -- successors 1406 
    -- members (6) 
      -- 	branch_block_stmt_2042/assign_stmt_2355_to_assign_stmt_2367__exit__
      -- 	branch_block_stmt_2042/bb_14_bbx_xnph7x_xix_xix_xi33
      -- 	branch_block_stmt_2042/assign_stmt_2355_to_assign_stmt_2367/OR_u32_u32_2366_Update/ca
      -- 	branch_block_stmt_2042/assign_stmt_2355_to_assign_stmt_2367/OR_u32_u32_2366_Update/$exit
      -- 	branch_block_stmt_2042/assign_stmt_2355_to_assign_stmt_2367/$exit
      -- 	branch_block_stmt_2042/assign_stmt_2355_to_assign_stmt_2367/OR_u32_u32_2366_update_completed_
      -- 
    ca_11472_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => OR_u32_u32_2366_inst_ack_1, ack => cp_elements(290)); -- 
    -- CP-element group 291 fork  transition  bypass 
    -- predecessors 12 
    -- successors 292 293 296 
    -- members (1) 
      -- 	branch_block_stmt_2042/assign_stmt_2389_to_assign_stmt_2395/$entry
      -- 
    cp_elements(291) <= cp_elements(12);
    -- CP-element group 292 transition  output  bypass 
    -- predecessors 291 
    -- successors 295 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_2389_to_assign_stmt_2395/LSHR_u32_u32_2388_Update/cr
      -- 	branch_block_stmt_2042/assign_stmt_2389_to_assign_stmt_2395/LSHR_u32_u32_2388_Update/$entry
      -- 	branch_block_stmt_2042/assign_stmt_2389_to_assign_stmt_2395/LSHR_u32_u32_2388_update_start_
      -- 
    cp_elements(292) <= cp_elements(291);
    cr_11492_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(292), ack => LSHR_u32_u32_2388_inst_req_1); -- 
    -- CP-element group 293 transition  output  bypass 
    -- predecessors 291 
    -- successors 294 
    -- members (7) 
      -- 	branch_block_stmt_2042/assign_stmt_2389_to_assign_stmt_2395/LSHR_u32_u32_2388_Sample/rr
      -- 	branch_block_stmt_2042/assign_stmt_2389_to_assign_stmt_2395/LSHR_u32_u32_2388_Sample/$entry
      -- 	branch_block_stmt_2042/assign_stmt_2389_to_assign_stmt_2395/R_xx_x016x_xix_xix_xi31_2385_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2389_to_assign_stmt_2395/R_xx_x016x_xix_xix_xi31_2385_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_2389_to_assign_stmt_2395/R_xx_x016x_xix_xix_xi31_2385_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2389_to_assign_stmt_2395/R_xx_x016x_xix_xix_xi31_2385_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_2389_to_assign_stmt_2395/LSHR_u32_u32_2388_sample_start_
      -- 
    cp_elements(293) <= cp_elements(291);
    rr_11487_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(293), ack => LSHR_u32_u32_2388_inst_req_0); -- 
    -- CP-element group 294 transition  input  bypass 
    -- predecessors 293 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_2389_to_assign_stmt_2395/LSHR_u32_u32_2388_Sample/ra
      -- 	branch_block_stmt_2042/assign_stmt_2389_to_assign_stmt_2395/LSHR_u32_u32_2388_Sample/$exit
      -- 	branch_block_stmt_2042/assign_stmt_2389_to_assign_stmt_2395/LSHR_u32_u32_2388_sample_completed_
      -- 
    ra_11488_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => LSHR_u32_u32_2388_inst_ack_0, ack => cp_elements(294)); -- 
    -- CP-element group 295 transition  input  output  bypass 
    -- predecessors 292 
    -- successors 297 
    -- members (10) 
      -- 	branch_block_stmt_2042/assign_stmt_2389_to_assign_stmt_2395/UGT_u32_u1_2394_Sample/$entry
      -- 	branch_block_stmt_2042/assign_stmt_2389_to_assign_stmt_2395/R_iNsTr_78_2391_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2389_to_assign_stmt_2395/R_iNsTr_78_2391_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_2389_to_assign_stmt_2395/UGT_u32_u1_2394_Sample/rr
      -- 	branch_block_stmt_2042/assign_stmt_2389_to_assign_stmt_2395/R_iNsTr_78_2391_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2389_to_assign_stmt_2395/R_iNsTr_78_2391_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_2389_to_assign_stmt_2395/UGT_u32_u1_2394_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_2389_to_assign_stmt_2395/LSHR_u32_u32_2388_Update/ca
      -- 	branch_block_stmt_2042/assign_stmt_2389_to_assign_stmt_2395/LSHR_u32_u32_2388_Update/$exit
      -- 	branch_block_stmt_2042/assign_stmt_2389_to_assign_stmt_2395/LSHR_u32_u32_2388_update_completed_
      -- 
    ca_11493_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => LSHR_u32_u32_2388_inst_ack_1, ack => cp_elements(295)); -- 
    rr_11505_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(295), ack => UGT_u32_u1_2394_inst_req_0); -- 
    -- CP-element group 296 transition  output  bypass 
    -- predecessors 291 
    -- successors 298 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_2389_to_assign_stmt_2395/UGT_u32_u1_2394_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_2389_to_assign_stmt_2395/UGT_u32_u1_2394_Update/$entry
      -- 	branch_block_stmt_2042/assign_stmt_2389_to_assign_stmt_2395/UGT_u32_u1_2394_Update/cr
      -- 
    cp_elements(296) <= cp_elements(291);
    cr_11510_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(296), ack => UGT_u32_u1_2394_inst_req_1); -- 
    -- CP-element group 297 transition  input  bypass 
    -- predecessors 295 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_2389_to_assign_stmt_2395/UGT_u32_u1_2394_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2389_to_assign_stmt_2395/UGT_u32_u1_2394_Sample/$exit
      -- 	branch_block_stmt_2042/assign_stmt_2389_to_assign_stmt_2395/UGT_u32_u1_2394_Sample/ra
      -- 
    ra_11506_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => UGT_u32_u1_2394_inst_ack_0, ack => cp_elements(297)); -- 
    -- CP-element group 298 branch  transition  place  input  bypass 
    -- predecessors 296 
    -- successors 299 300 
    -- members (6) 
      -- 	branch_block_stmt_2042/assign_stmt_2389_to_assign_stmt_2395/UGT_u32_u1_2394_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2389_to_assign_stmt_2395/UGT_u32_u1_2394_Update/$exit
      -- 	branch_block_stmt_2042/assign_stmt_2389_to_assign_stmt_2395/UGT_u32_u1_2394_Update/ca
      -- 	branch_block_stmt_2042/assign_stmt_2389_to_assign_stmt_2395__exit__
      -- 	branch_block_stmt_2042/if_stmt_2396__entry__
      -- 	branch_block_stmt_2042/assign_stmt_2389_to_assign_stmt_2395/$exit
      -- 
    ca_11511_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => UGT_u32_u1_2394_inst_ack_1, ack => cp_elements(298)); -- 
    -- CP-element group 299 transition  place  dead  bypass 
    -- predecessors 298 
    -- successors 13 
    -- members (8) 
      -- 	branch_block_stmt_2042/if_stmt_2396_dead_link/$entry
      -- 	branch_block_stmt_2042/if_stmt_2396_dead_link/$exit
      -- 	branch_block_stmt_2042/if_stmt_2396_dead_link/dead_transition
      -- 	branch_block_stmt_2042/if_stmt_2396__exit__
      -- 	branch_block_stmt_2042/merge_stmt_2402__entry__
      -- 	branch_block_stmt_2042/merge_stmt_2402_dead_link/$entry
      -- 	branch_block_stmt_2042/merge_stmt_2402_dead_link/$exit
      -- 	branch_block_stmt_2042/merge_stmt_2402_dead_link/dead_transition
      -- 
    cp_elements(299) <= false;
    -- CP-element group 300 transition  output  bypass 
    -- predecessors 298 
    -- successors 301 
    -- members (3) 
      -- 	branch_block_stmt_2042/if_stmt_2396_eval_test/$entry
      -- 	branch_block_stmt_2042/if_stmt_2396_eval_test/$exit
      -- 	branch_block_stmt_2042/if_stmt_2396_eval_test/branch_req
      -- 
    cp_elements(300) <= cp_elements(298);
    branch_req_11519_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(300), ack => if_stmt_2396_branch_req_0); -- 
    -- CP-element group 301 branch  place  bypass 
    -- predecessors 300 
    -- successors 302 304 
    -- members (1) 
      -- 	branch_block_stmt_2042/R_iNsTr_79_2397_place
      -- 
    cp_elements(301) <= cp_elements(300);
    -- CP-element group 302 transition  bypass 
    -- predecessors 301 
    -- successors 303 
    -- members (1) 
      -- 	branch_block_stmt_2042/if_stmt_2396_if_link/$entry
      -- 
    cp_elements(302) <= cp_elements(301);
    -- CP-element group 303 transition  place  input  bypass 
    -- predecessors 302 
    -- successors 13 
    -- members (9) 
      -- 	branch_block_stmt_2042/if_stmt_2396_if_link/$exit
      -- 	branch_block_stmt_2042/if_stmt_2396_if_link/if_choice_transition
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xix_xi33_bbx_xnphx_xix_xix_xi36x_xpreheader
      -- 	branch_block_stmt_2042/merge_stmt_2402_PhiReqMerge
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xix_xi33_bbx_xnphx_xix_xix_xi36x_xpreheader_PhiReq/$entry
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xix_xi33_bbx_xnphx_xix_xix_xi36x_xpreheader_PhiReq/$exit
      -- 	branch_block_stmt_2042/merge_stmt_2402_PhiAck/$entry
      -- 	branch_block_stmt_2042/merge_stmt_2402_PhiAck/$exit
      -- 	branch_block_stmt_2042/merge_stmt_2402_PhiAck/dummy
      -- 
    if_choice_transition_11524_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2396_branch_ack_1, ack => cp_elements(303)); -- 
    -- CP-element group 304 transition  bypass 
    -- predecessors 301 
    -- successors 305 
    -- members (1) 
      -- 	branch_block_stmt_2042/if_stmt_2396_else_link/$entry
      -- 
    cp_elements(304) <= cp_elements(301);
    -- CP-element group 305 transition  place  input  bypass 
    -- predecessors 304 
    -- successors 1497 
    -- members (3) 
      -- 	branch_block_stmt_2042/if_stmt_2396_else_link/$exit
      -- 	branch_block_stmt_2042/if_stmt_2396_else_link/else_choice_transition
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xix_xi33_xx_x_crit_edgex_xix_xix_xi39
      -- 
    else_choice_transition_11528_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2396_branch_ack_0, ack => cp_elements(305)); -- 
    -- CP-element group 306 fork  transition  bypass 
    -- predecessors 14 
    -- successors 307 308 311 312 316 317 
    -- members (1) 
      -- 	branch_block_stmt_2042/assign_stmt_2425_to_assign_stmt_2436/$entry
      -- 
    cp_elements(306) <= cp_elements(14);
    -- CP-element group 307 transition  output  bypass 
    -- predecessors 306 
    -- successors 310 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_2425_to_assign_stmt_2436/SHL_u32_u32_2424_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_2425_to_assign_stmt_2436/SHL_u32_u32_2424_Update/$entry
      -- 	branch_block_stmt_2042/assign_stmt_2425_to_assign_stmt_2436/SHL_u32_u32_2424_Update/cr
      -- 
    cp_elements(307) <= cp_elements(306);
    cr_11550_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(307), ack => SHL_u32_u32_2424_inst_req_1); -- 
    -- CP-element group 308 transition  output  bypass 
    -- predecessors 306 
    -- successors 309 
    -- members (7) 
      -- 	branch_block_stmt_2042/assign_stmt_2425_to_assign_stmt_2436/SHL_u32_u32_2424_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_2425_to_assign_stmt_2436/R_shifted_divisorx_x03x_xix_xix_xi34_2421_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_2425_to_assign_stmt_2436/R_shifted_divisorx_x03x_xix_xix_xi34_2421_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2425_to_assign_stmt_2436/R_shifted_divisorx_x03x_xix_xix_xi34_2421_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_2425_to_assign_stmt_2436/R_shifted_divisorx_x03x_xix_xix_xi34_2421_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2425_to_assign_stmt_2436/SHL_u32_u32_2424_Sample/$entry
      -- 	branch_block_stmt_2042/assign_stmt_2425_to_assign_stmt_2436/SHL_u32_u32_2424_Sample/rr
      -- 
    cp_elements(308) <= cp_elements(306);
    rr_11545_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(308), ack => SHL_u32_u32_2424_inst_req_0); -- 
    -- CP-element group 309 transition  input  bypass 
    -- predecessors 308 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_2425_to_assign_stmt_2436/SHL_u32_u32_2424_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2425_to_assign_stmt_2436/SHL_u32_u32_2424_Sample/$exit
      -- 	branch_block_stmt_2042/assign_stmt_2425_to_assign_stmt_2436/SHL_u32_u32_2424_Sample/ra
      -- 
    ra_11546_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => SHL_u32_u32_2424_inst_ack_0, ack => cp_elements(309)); -- 
    -- CP-element group 310 transition  input  bypass 
    -- predecessors 307 
    -- successors 315 
    -- members (7) 
      -- 	branch_block_stmt_2042/assign_stmt_2425_to_assign_stmt_2436/SHL_u32_u32_2424_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2425_to_assign_stmt_2436/SHL_u32_u32_2424_Update/$exit
      -- 	branch_block_stmt_2042/assign_stmt_2425_to_assign_stmt_2436/R_iNsTr_135_2433_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2425_to_assign_stmt_2436/R_iNsTr_135_2433_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_2425_to_assign_stmt_2436/R_iNsTr_135_2433_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2425_to_assign_stmt_2436/R_iNsTr_135_2433_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_2425_to_assign_stmt_2436/SHL_u32_u32_2424_Update/ca
      -- 
    ca_11551_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => SHL_u32_u32_2424_inst_ack_1, ack => cp_elements(310)); -- 
    -- CP-element group 311 transition  output  bypass 
    -- predecessors 306 
    -- successors 314 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_2425_to_assign_stmt_2436/SHL_u32_u32_2430_Update/$entry
      -- 	branch_block_stmt_2042/assign_stmt_2425_to_assign_stmt_2436/SHL_u32_u32_2430_Update/cr
      -- 	branch_block_stmt_2042/assign_stmt_2425_to_assign_stmt_2436/SHL_u32_u32_2430_update_start_
      -- 
    cp_elements(311) <= cp_elements(306);
    cr_11568_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(311), ack => SHL_u32_u32_2430_inst_req_1); -- 
    -- CP-element group 312 transition  output  bypass 
    -- predecessors 306 
    -- successors 313 
    -- members (7) 
      -- 	branch_block_stmt_2042/assign_stmt_2425_to_assign_stmt_2436/SHL_u32_u32_2430_Sample/$entry
      -- 	branch_block_stmt_2042/assign_stmt_2425_to_assign_stmt_2436/R_curr_quotientx_x02x_xix_xix_xi35_2427_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2425_to_assign_stmt_2436/R_curr_quotientx_x02x_xix_xix_xi35_2427_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_2425_to_assign_stmt_2436/SHL_u32_u32_2430_Sample/rr
      -- 	branch_block_stmt_2042/assign_stmt_2425_to_assign_stmt_2436/R_curr_quotientx_x02x_xix_xix_xi35_2427_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2425_to_assign_stmt_2436/R_curr_quotientx_x02x_xix_xix_xi35_2427_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_2425_to_assign_stmt_2436/SHL_u32_u32_2430_sample_start_
      -- 
    cp_elements(312) <= cp_elements(306);
    rr_11563_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(312), ack => SHL_u32_u32_2430_inst_req_0); -- 
    -- CP-element group 313 transition  input  bypass 
    -- predecessors 312 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_2425_to_assign_stmt_2436/SHL_u32_u32_2430_Sample/$exit
      -- 	branch_block_stmt_2042/assign_stmt_2425_to_assign_stmt_2436/SHL_u32_u32_2430_Sample/ra
      -- 	branch_block_stmt_2042/assign_stmt_2425_to_assign_stmt_2436/SHL_u32_u32_2430_sample_completed_
      -- 
    ra_11564_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => SHL_u32_u32_2430_inst_ack_0, ack => cp_elements(313)); -- 
    -- CP-element group 314 transition  input  bypass 
    -- predecessors 311 
    -- successors 320 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_2425_to_assign_stmt_2436/SHL_u32_u32_2430_Update/$exit
      -- 	branch_block_stmt_2042/assign_stmt_2425_to_assign_stmt_2436/SHL_u32_u32_2430_Update/ca
      -- 	branch_block_stmt_2042/assign_stmt_2425_to_assign_stmt_2436/SHL_u32_u32_2430_update_completed_
      -- 
    ca_11569_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => SHL_u32_u32_2430_inst_ack_1, ack => cp_elements(314)); -- 
    -- CP-element group 315 join  transition  output  bypass 
    -- predecessors 310 317 
    -- successors 318 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_2425_to_assign_stmt_2436/ULT_u32_u1_2435_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_2425_to_assign_stmt_2436/ULT_u32_u1_2435_Sample/rr
      -- 	branch_block_stmt_2042/assign_stmt_2425_to_assign_stmt_2436/ULT_u32_u1_2435_Sample/$entry
      -- 
    cp_element_group_315: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 20) := "cp_element_group_315"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(310) & cp_elements(317);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(315), clk => clk, reset => reset); --
    end block;
    rr_11585_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(315), ack => ULT_u32_u1_2435_inst_req_0); -- 
    -- CP-element group 316 transition  output  bypass 
    -- predecessors 306 
    -- successors 319 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_2425_to_assign_stmt_2436/ULT_u32_u1_2435_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_2425_to_assign_stmt_2436/ULT_u32_u1_2435_Update/$entry
      -- 	branch_block_stmt_2042/assign_stmt_2425_to_assign_stmt_2436/ULT_u32_u1_2435_Update/cr
      -- 
    cp_elements(316) <= cp_elements(306);
    cr_11590_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(316), ack => ULT_u32_u1_2435_inst_req_1); -- 
    -- CP-element group 317 transition  bypass 
    -- predecessors 306 
    -- successors 315 
    -- members (4) 
      -- 	branch_block_stmt_2042/assign_stmt_2425_to_assign_stmt_2436/R_iNsTr_78_2434_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_2425_to_assign_stmt_2436/R_iNsTr_78_2434_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2425_to_assign_stmt_2436/R_iNsTr_78_2434_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_2425_to_assign_stmt_2436/R_iNsTr_78_2434_sample_completed_
      -- 
    cp_elements(317) <= cp_elements(306);
    -- CP-element group 318 transition  input  bypass 
    -- predecessors 315 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_2425_to_assign_stmt_2436/ULT_u32_u1_2435_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2425_to_assign_stmt_2436/ULT_u32_u1_2435_Sample/ra
      -- 	branch_block_stmt_2042/assign_stmt_2425_to_assign_stmt_2436/ULT_u32_u1_2435_Sample/$exit
      -- 
    ra_11586_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ULT_u32_u1_2435_inst_ack_0, ack => cp_elements(318)); -- 
    -- CP-element group 319 transition  input  bypass 
    -- predecessors 316 
    -- successors 320 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_2425_to_assign_stmt_2436/ULT_u32_u1_2435_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2425_to_assign_stmt_2436/ULT_u32_u1_2435_Update/ca
      -- 	branch_block_stmt_2042/assign_stmt_2425_to_assign_stmt_2436/ULT_u32_u1_2435_Update/$exit
      -- 
    ca_11591_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ULT_u32_u1_2435_inst_ack_1, ack => cp_elements(319)); -- 
    -- CP-element group 320 join  transition  bypass 
    -- predecessors 314 319 
    -- successors 15 
    -- members (1) 
      -- 	branch_block_stmt_2042/assign_stmt_2425_to_assign_stmt_2436/$exit
      -- 
    cp_element_group_320: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 20) := "cp_element_group_320"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(314) & cp_elements(319);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(320), clk => clk, reset => reset); --
    end block;
    -- CP-element group 321 transition  place  dead  bypass 
    -- predecessors 15 
    -- successors 16 
    -- members (8) 
      -- 	branch_block_stmt_2042/if_stmt_2437__exit__
      -- 	branch_block_stmt_2042/merge_stmt_2443__entry__
      -- 	branch_block_stmt_2042/if_stmt_2437_dead_link/dead_transition
      -- 	branch_block_stmt_2042/if_stmt_2437_dead_link/$exit
      -- 	branch_block_stmt_2042/if_stmt_2437_dead_link/$entry
      -- 	branch_block_stmt_2042/merge_stmt_2443_dead_link/$entry
      -- 	branch_block_stmt_2042/merge_stmt_2443_dead_link/$exit
      -- 	branch_block_stmt_2042/merge_stmt_2443_dead_link/dead_transition
      -- 
    cp_elements(321) <= false;
    -- CP-element group 322 transition  output  bypass 
    -- predecessors 15 
    -- successors 323 
    -- members (3) 
      -- 	branch_block_stmt_2042/if_stmt_2437_eval_test/$exit
      -- 	branch_block_stmt_2042/if_stmt_2437_eval_test/branch_req
      -- 	branch_block_stmt_2042/if_stmt_2437_eval_test/$entry
      -- 
    cp_elements(322) <= cp_elements(15);
    branch_req_11599_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(322), ack => if_stmt_2437_branch_req_0); -- 
    -- CP-element group 323 branch  place  bypass 
    -- predecessors 322 
    -- successors 324 326 
    -- members (1) 
      -- 	branch_block_stmt_2042/R_iNsTr_137_2438_place
      -- 
    cp_elements(323) <= cp_elements(322);
    -- CP-element group 324 transition  bypass 
    -- predecessors 323 
    -- successors 325 
    -- members (1) 
      -- 	branch_block_stmt_2042/if_stmt_2437_if_link/$entry
      -- 
    cp_elements(324) <= cp_elements(323);
    -- CP-element group 325 transition  place  input  bypass 
    -- predecessors 324 
    -- successors 1449 
    -- members (3) 
      -- 	branch_block_stmt_2042/if_stmt_2437_if_link/if_choice_transition
      -- 	branch_block_stmt_2042/if_stmt_2437_if_link/$exit
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi36_bbx_xnphx_xix_xix_xi36
      -- 
    if_choice_transition_11604_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2437_branch_ack_1, ack => cp_elements(325)); -- 
    -- CP-element group 326 transition  bypass 
    -- predecessors 323 
    -- successors 327 
    -- members (1) 
      -- 	branch_block_stmt_2042/if_stmt_2437_else_link/$entry
      -- 
    cp_elements(326) <= cp_elements(323);
    -- CP-element group 327 transition  place  input  bypass 
    -- predecessors 326 
    -- successors 1478 
    -- members (3) 
      -- 	branch_block_stmt_2042/if_stmt_2437_else_link/$exit
      -- 	branch_block_stmt_2042/if_stmt_2437_else_link/else_choice_transition
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi36_xx_x_crit_edgex_xix_xix_xi39x_xloopexit
      -- 
    else_choice_transition_11608_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2437_branch_ack_0, ack => cp_elements(327)); -- 
    -- CP-element group 328 fork  transition  bypass 
    -- predecessors 17 
    -- successors 330 331 332 336 337 338 341 
    -- members (1) 
      -- 	branch_block_stmt_2042/assign_stmt_2474_to_assign_stmt_2485/$entry
      -- 
    cp_elements(328) <= cp_elements(17);
    -- CP-element group 329 join  transition  output  bypass 
    -- predecessors 331 332 
    -- successors 333 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_2474_to_assign_stmt_2485/ADD_u32_u32_2473_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_2474_to_assign_stmt_2485/ADD_u32_u32_2473_Sample/$entry
      -- 	branch_block_stmt_2042/assign_stmt_2474_to_assign_stmt_2485/ADD_u32_u32_2473_Sample/rr
      -- 
    cp_element_group_329: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 20) := "cp_element_group_329"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(331) & cp_elements(332);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(329), clk => clk, reset => reset); --
    end block;
    rr_11629_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(329), ack => ADD_u32_u32_2473_inst_req_0); -- 
    -- CP-element group 330 transition  output  bypass 
    -- predecessors 328 
    -- successors 334 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_2474_to_assign_stmt_2485/ADD_u32_u32_2473_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_2474_to_assign_stmt_2485/ADD_u32_u32_2473_Update/$entry
      -- 	branch_block_stmt_2042/assign_stmt_2474_to_assign_stmt_2485/ADD_u32_u32_2473_Update/cr
      -- 
    cp_elements(330) <= cp_elements(328);
    cr_11634_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(330), ack => ADD_u32_u32_2473_inst_req_1); -- 
    -- CP-element group 331 transition  bypass 
    -- predecessors 328 
    -- successors 329 
    -- members (4) 
      -- 	branch_block_stmt_2042/assign_stmt_2474_to_assign_stmt_2485/R_curr_quotientx_x0x_xlcssax_xix_xix_xi38_2471_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2474_to_assign_stmt_2485/R_curr_quotientx_x0x_xlcssax_xix_xix_xi38_2471_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2474_to_assign_stmt_2485/R_curr_quotientx_x0x_xlcssax_xix_xix_xi38_2471_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_2474_to_assign_stmt_2485/R_curr_quotientx_x0x_xlcssax_xix_xix_xi38_2471_sample_start_
      -- 
    cp_elements(331) <= cp_elements(328);
    -- CP-element group 332 transition  bypass 
    -- predecessors 328 
    -- successors 329 
    -- members (4) 
      -- 	branch_block_stmt_2042/assign_stmt_2474_to_assign_stmt_2485/R_quotientx_x05x_xix_xix_xi32_2472_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_2474_to_assign_stmt_2485/R_quotientx_x05x_xix_xix_xi32_2472_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2474_to_assign_stmt_2485/R_quotientx_x05x_xix_xix_xi32_2472_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_2474_to_assign_stmt_2485/R_quotientx_x05x_xix_xix_xi32_2472_sample_completed_
      -- 
    cp_elements(332) <= cp_elements(328);
    -- CP-element group 333 transition  input  bypass 
    -- predecessors 329 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_2474_to_assign_stmt_2485/ADD_u32_u32_2473_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2474_to_assign_stmt_2485/ADD_u32_u32_2473_Sample/$exit
      -- 	branch_block_stmt_2042/assign_stmt_2474_to_assign_stmt_2485/ADD_u32_u32_2473_Sample/ra
      -- 
    ra_11630_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u32_u32_2473_inst_ack_0, ack => cp_elements(333)); -- 
    -- CP-element group 334 transition  input  bypass 
    -- predecessors 330 
    -- successors 344 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_2474_to_assign_stmt_2485/ADD_u32_u32_2473_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2474_to_assign_stmt_2485/ADD_u32_u32_2473_Update/$exit
      -- 	branch_block_stmt_2042/assign_stmt_2474_to_assign_stmt_2485/ADD_u32_u32_2473_Update/ca
      -- 
    ca_11635_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u32_u32_2473_inst_ack_1, ack => cp_elements(334)); -- 
    -- CP-element group 335 join  transition  output  bypass 
    -- predecessors 337 338 
    -- successors 339 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_2474_to_assign_stmt_2485/SUB_u32_u32_2478_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_2474_to_assign_stmt_2485/SUB_u32_u32_2478_Sample/$entry
      -- 	branch_block_stmt_2042/assign_stmt_2474_to_assign_stmt_2485/SUB_u32_u32_2478_Sample/rr
      -- 
    cp_element_group_335: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 20) := "cp_element_group_335"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(337) & cp_elements(338);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(335), clk => clk, reset => reset); --
    end block;
    rr_11651_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(335), ack => SUB_u32_u32_2478_inst_req_0); -- 
    -- CP-element group 336 transition  output  bypass 
    -- predecessors 328 
    -- successors 340 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_2474_to_assign_stmt_2485/SUB_u32_u32_2478_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_2474_to_assign_stmt_2485/SUB_u32_u32_2478_Update/$entry
      -- 	branch_block_stmt_2042/assign_stmt_2474_to_assign_stmt_2485/SUB_u32_u32_2478_Update/cr
      -- 
    cp_elements(336) <= cp_elements(328);
    cr_11656_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(336), ack => SUB_u32_u32_2478_inst_req_1); -- 
    -- CP-element group 337 transition  bypass 
    -- predecessors 328 
    -- successors 335 
    -- members (4) 
      -- 	branch_block_stmt_2042/assign_stmt_2474_to_assign_stmt_2485/R_xx_x016x_xix_xix_xi31_2476_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_2474_to_assign_stmt_2485/R_xx_x016x_xix_xix_xi31_2476_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2474_to_assign_stmt_2485/R_xx_x016x_xix_xix_xi31_2476_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_2474_to_assign_stmt_2485/R_xx_x016x_xix_xix_xi31_2476_update_completed_
      -- 
    cp_elements(337) <= cp_elements(328);
    -- CP-element group 338 transition  bypass 
    -- predecessors 328 
    -- successors 335 
    -- members (4) 
      -- 	branch_block_stmt_2042/assign_stmt_2474_to_assign_stmt_2485/R_shifted_divisorx_x0x_xlcssax_xix_xix_xi37_2477_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_2474_to_assign_stmt_2485/R_shifted_divisorx_x0x_xlcssax_xix_xix_xi37_2477_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2474_to_assign_stmt_2485/R_shifted_divisorx_x0x_xlcssax_xix_xix_xi37_2477_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_2474_to_assign_stmt_2485/R_shifted_divisorx_x0x_xlcssax_xix_xix_xi37_2477_update_completed_
      -- 
    cp_elements(338) <= cp_elements(328);
    -- CP-element group 339 transition  input  bypass 
    -- predecessors 335 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_2474_to_assign_stmt_2485/SUB_u32_u32_2478_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2474_to_assign_stmt_2485/SUB_u32_u32_2478_Sample/$exit
      -- 	branch_block_stmt_2042/assign_stmt_2474_to_assign_stmt_2485/SUB_u32_u32_2478_Sample/ra
      -- 
    ra_11652_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => SUB_u32_u32_2478_inst_ack_0, ack => cp_elements(339)); -- 
    -- CP-element group 340 transition  input  output  bypass 
    -- predecessors 336 
    -- successors 342 
    -- members (10) 
      -- 	branch_block_stmt_2042/assign_stmt_2474_to_assign_stmt_2485/SUB_u32_u32_2478_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2474_to_assign_stmt_2485/SUB_u32_u32_2478_Update/$exit
      -- 	branch_block_stmt_2042/assign_stmt_2474_to_assign_stmt_2485/SUB_u32_u32_2478_Update/ca
      -- 	branch_block_stmt_2042/assign_stmt_2474_to_assign_stmt_2485/ULT_u32_u1_2484_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_2474_to_assign_stmt_2485/R_iNsTr_110_2481_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_2474_to_assign_stmt_2485/R_iNsTr_110_2481_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2474_to_assign_stmt_2485/R_iNsTr_110_2481_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_2474_to_assign_stmt_2485/R_iNsTr_110_2481_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2474_to_assign_stmt_2485/ULT_u32_u1_2484_Sample/$entry
      -- 	branch_block_stmt_2042/assign_stmt_2474_to_assign_stmt_2485/ULT_u32_u1_2484_Sample/rr
      -- 
    ca_11657_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => SUB_u32_u32_2478_inst_ack_1, ack => cp_elements(340)); -- 
    rr_11669_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(340), ack => ULT_u32_u1_2484_inst_req_0); -- 
    -- CP-element group 341 transition  output  bypass 
    -- predecessors 328 
    -- successors 343 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_2474_to_assign_stmt_2485/ULT_u32_u1_2484_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_2474_to_assign_stmt_2485/ULT_u32_u1_2484_Update/$entry
      -- 	branch_block_stmt_2042/assign_stmt_2474_to_assign_stmt_2485/ULT_u32_u1_2484_Update/cr
      -- 
    cp_elements(341) <= cp_elements(328);
    cr_11674_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(341), ack => ULT_u32_u1_2484_inst_req_1); -- 
    -- CP-element group 342 transition  input  bypass 
    -- predecessors 340 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_2474_to_assign_stmt_2485/ULT_u32_u1_2484_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2474_to_assign_stmt_2485/ULT_u32_u1_2484_Sample/$exit
      -- 	branch_block_stmt_2042/assign_stmt_2474_to_assign_stmt_2485/ULT_u32_u1_2484_Sample/ra
      -- 
    ra_11670_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ULT_u32_u1_2484_inst_ack_0, ack => cp_elements(342)); -- 
    -- CP-element group 343 transition  input  bypass 
    -- predecessors 341 
    -- successors 344 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_2474_to_assign_stmt_2485/ULT_u32_u1_2484_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2474_to_assign_stmt_2485/ULT_u32_u1_2484_Update/$exit
      -- 	branch_block_stmt_2042/assign_stmt_2474_to_assign_stmt_2485/ULT_u32_u1_2484_Update/ca
      -- 
    ca_11675_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ULT_u32_u1_2484_inst_ack_1, ack => cp_elements(343)); -- 
    -- CP-element group 344 join  transition  bypass 
    -- predecessors 334 343 
    -- successors 18 
    -- members (1) 
      -- 	branch_block_stmt_2042/assign_stmt_2474_to_assign_stmt_2485/$exit
      -- 
    cp_element_group_344: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 20) := "cp_element_group_344"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(334) & cp_elements(343);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(344), clk => clk, reset => reset); --
    end block;
    -- CP-element group 345 transition  place  dead  bypass 
    -- predecessors 18 
    -- successors 19 
    -- members (8) 
      -- 	branch_block_stmt_2042/if_stmt_2486__exit__
      -- 	branch_block_stmt_2042/merge_stmt_2492__entry__
      -- 	branch_block_stmt_2042/if_stmt_2486_dead_link/$entry
      -- 	branch_block_stmt_2042/if_stmt_2486_dead_link/$exit
      -- 	branch_block_stmt_2042/if_stmt_2486_dead_link/dead_transition
      -- 	branch_block_stmt_2042/merge_stmt_2492_dead_link/$entry
      -- 	branch_block_stmt_2042/merge_stmt_2492_dead_link/$exit
      -- 	branch_block_stmt_2042/merge_stmt_2492_dead_link/dead_transition
      -- 
    cp_elements(345) <= false;
    -- CP-element group 346 transition  output  bypass 
    -- predecessors 18 
    -- successors 347 
    -- members (3) 
      -- 	branch_block_stmt_2042/if_stmt_2486_eval_test/$entry
      -- 	branch_block_stmt_2042/if_stmt_2486_eval_test/$exit
      -- 	branch_block_stmt_2042/if_stmt_2486_eval_test/branch_req
      -- 
    cp_elements(346) <= cp_elements(18);
    branch_req_11683_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(346), ack => if_stmt_2486_branch_req_0); -- 
    -- CP-element group 347 branch  place  bypass 
    -- predecessors 346 
    -- successors 348 350 
    -- members (1) 
      -- 	branch_block_stmt_2042/R_iNsTr_111_2487_place
      -- 
    cp_elements(347) <= cp_elements(346);
    -- CP-element group 348 transition  bypass 
    -- predecessors 347 
    -- successors 349 
    -- members (1) 
      -- 	branch_block_stmt_2042/if_stmt_2486_if_link/$entry
      -- 
    cp_elements(348) <= cp_elements(347);
    -- CP-element group 349 fork  transition  place  input  bypass 
    -- predecessors 348 
    -- successors 1526 1528 
    -- members (8) 
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi39_udiv32x_xexitx_xpreheaderx_xix_xi41
      -- 	branch_block_stmt_2042/if_stmt_2486_if_link/$exit
      -- 	branch_block_stmt_2042/if_stmt_2486_if_link/if_choice_transition
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi39_udiv32x_xexitx_xpreheaderx_xix_xi41_PhiReq/$entry
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi39_udiv32x_xexitx_xpreheaderx_xix_xi41_PhiReq/phi_stmt_2493/$entry
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi39_udiv32x_xexitx_xpreheaderx_xix_xi41_PhiReq/phi_stmt_2493/phi_stmt_2493_sources/$entry
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi39_udiv32x_xexitx_xpreheaderx_xix_xi41_PhiReq/phi_stmt_2493/phi_stmt_2493_sources/type_cast_2496/$entry
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi39_udiv32x_xexitx_xpreheaderx_xix_xi41_PhiReq/phi_stmt_2493/phi_stmt_2493_sources/type_cast_2496/SplitProtocol/$entry
      -- 
    if_choice_transition_11688_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2486_branch_ack_1, ack => cp_elements(349)); -- 
    -- CP-element group 350 transition  bypass 
    -- predecessors 347 
    -- successors 351 
    -- members (1) 
      -- 	branch_block_stmt_2042/if_stmt_2486_else_link/$entry
      -- 
    cp_elements(350) <= cp_elements(347);
    -- CP-element group 351 transition  place  input  bypass 
    -- predecessors 350 
    -- successors 1424 
    -- members (3) 
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi39_bbx_xnph7x_xix_xix_xi33
      -- 	branch_block_stmt_2042/if_stmt_2486_else_link/$exit
      -- 	branch_block_stmt_2042/if_stmt_2486_else_link/else_choice_transition
      -- 
    else_choice_transition_11692_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2486_branch_ack_0, ack => cp_elements(351)); -- 
    -- CP-element group 352 fork  transition  bypass 
    -- predecessors 19 
    -- successors 353 354 357 358 361 364 367 368 371 374 375 381 
    -- members (1) 
      -- 	branch_block_stmt_2042/assign_stmt_2503_to_assign_stmt_2546/$entry
      -- 
    cp_elements(352) <= cp_elements(19);
    -- CP-element group 353 transition  output  bypass 
    -- predecessors 352 
    -- successors 356 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_2503_to_assign_stmt_2546/LSHR_u32_u32_2502_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_2503_to_assign_stmt_2546/LSHR_u32_u32_2502_Update/$entry
      -- 	branch_block_stmt_2042/assign_stmt_2503_to_assign_stmt_2546/LSHR_u32_u32_2502_Update/cr
      -- 
    cp_elements(353) <= cp_elements(352);
    cr_11714_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(353), ack => LSHR_u32_u32_2502_inst_req_1); -- 
    -- CP-element group 354 transition  output  bypass 
    -- predecessors 352 
    -- successors 355 
    -- members (7) 
      -- 	branch_block_stmt_2042/assign_stmt_2503_to_assign_stmt_2546/LSHR_u32_u32_2502_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_2503_to_assign_stmt_2546/R_tmp10x_xix_xi30_2499_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_2503_to_assign_stmt_2546/R_tmp10x_xix_xi30_2499_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2503_to_assign_stmt_2546/R_tmp10x_xix_xi30_2499_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_2503_to_assign_stmt_2546/R_tmp10x_xix_xi30_2499_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2503_to_assign_stmt_2546/LSHR_u32_u32_2502_Sample/$entry
      -- 	branch_block_stmt_2042/assign_stmt_2503_to_assign_stmt_2546/LSHR_u32_u32_2502_Sample/rr
      -- 
    cp_elements(354) <= cp_elements(352);
    rr_11709_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(354), ack => LSHR_u32_u32_2502_inst_req_0); -- 
    -- CP-element group 355 transition  input  bypass 
    -- predecessors 354 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_2503_to_assign_stmt_2546/LSHR_u32_u32_2502_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2503_to_assign_stmt_2546/LSHR_u32_u32_2502_Sample/$exit
      -- 	branch_block_stmt_2042/assign_stmt_2503_to_assign_stmt_2546/LSHR_u32_u32_2502_Sample/ra
      -- 
    ra_11710_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => LSHR_u32_u32_2502_inst_ack_0, ack => cp_elements(355)); -- 
    -- CP-element group 356 transition  input  output  bypass 
    -- predecessors 353 
    -- successors 362 
    -- members (10) 
      -- 	branch_block_stmt_2042/assign_stmt_2503_to_assign_stmt_2546/LSHR_u32_u32_2502_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2503_to_assign_stmt_2546/LSHR_u32_u32_2502_Update/$exit
      -- 	branch_block_stmt_2042/assign_stmt_2503_to_assign_stmt_2546/LSHR_u32_u32_2502_Update/ca
      -- 	branch_block_stmt_2042/assign_stmt_2503_to_assign_stmt_2546/AND_u32_u32_2514_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_2503_to_assign_stmt_2546/R_iNsTr_139_2511_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_2503_to_assign_stmt_2546/R_iNsTr_139_2511_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2503_to_assign_stmt_2546/R_iNsTr_139_2511_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_2503_to_assign_stmt_2546/R_iNsTr_139_2511_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2503_to_assign_stmt_2546/AND_u32_u32_2514_Sample/$entry
      -- 	branch_block_stmt_2042/assign_stmt_2503_to_assign_stmt_2546/AND_u32_u32_2514_Sample/rr
      -- 
    ca_11715_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => LSHR_u32_u32_2502_inst_ack_1, ack => cp_elements(356)); -- 
    rr_11745_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(356), ack => AND_u32_u32_2514_inst_req_0); -- 
    -- CP-element group 357 transition  output  bypass 
    -- predecessors 352 
    -- successors 360 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_2503_to_assign_stmt_2546/AND_u32_u32_2508_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_2503_to_assign_stmt_2546/AND_u32_u32_2508_Update/$entry
      -- 	branch_block_stmt_2042/assign_stmt_2503_to_assign_stmt_2546/AND_u32_u32_2508_Update/cr
      -- 
    cp_elements(357) <= cp_elements(352);
    cr_11732_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(357), ack => AND_u32_u32_2508_inst_req_1); -- 
    -- CP-element group 358 transition  output  bypass 
    -- predecessors 352 
    -- successors 359 
    -- members (7) 
      -- 	branch_block_stmt_2042/assign_stmt_2503_to_assign_stmt_2546/AND_u32_u32_2508_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_2503_to_assign_stmt_2546/R_tmp10x_xix_xi30_2505_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_2503_to_assign_stmt_2546/R_tmp10x_xix_xi30_2505_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2503_to_assign_stmt_2546/R_tmp10x_xix_xi30_2505_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_2503_to_assign_stmt_2546/R_tmp10x_xix_xi30_2505_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2503_to_assign_stmt_2546/AND_u32_u32_2508_Sample/$entry
      -- 	branch_block_stmt_2042/assign_stmt_2503_to_assign_stmt_2546/AND_u32_u32_2508_Sample/rr
      -- 
    cp_elements(358) <= cp_elements(352);
    rr_11727_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(358), ack => AND_u32_u32_2508_inst_req_0); -- 
    -- CP-element group 359 transition  input  bypass 
    -- predecessors 358 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_2503_to_assign_stmt_2546/AND_u32_u32_2508_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2503_to_assign_stmt_2546/AND_u32_u32_2508_Sample/$exit
      -- 	branch_block_stmt_2042/assign_stmt_2503_to_assign_stmt_2546/AND_u32_u32_2508_Sample/ra
      -- 
    ra_11728_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => AND_u32_u32_2508_inst_ack_0, ack => cp_elements(359)); -- 
    -- CP-element group 360 transition  input  bypass 
    -- predecessors 357 
    -- successors 384 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_2503_to_assign_stmt_2546/AND_u32_u32_2508_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2503_to_assign_stmt_2546/AND_u32_u32_2508_Update/$exit
      -- 	branch_block_stmt_2042/assign_stmt_2503_to_assign_stmt_2546/AND_u32_u32_2508_Update/ca
      -- 
    ca_11733_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => AND_u32_u32_2508_inst_ack_1, ack => cp_elements(360)); -- 
    -- CP-element group 361 transition  output  bypass 
    -- predecessors 352 
    -- successors 363 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_2503_to_assign_stmt_2546/AND_u32_u32_2514_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_2503_to_assign_stmt_2546/AND_u32_u32_2514_Update/$entry
      -- 	branch_block_stmt_2042/assign_stmt_2503_to_assign_stmt_2546/AND_u32_u32_2514_Update/cr
      -- 
    cp_elements(361) <= cp_elements(352);
    cr_11750_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(361), ack => AND_u32_u32_2514_inst_req_1); -- 
    -- CP-element group 362 transition  input  bypass 
    -- predecessors 356 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_2503_to_assign_stmt_2546/AND_u32_u32_2514_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2503_to_assign_stmt_2546/AND_u32_u32_2514_Sample/$exit
      -- 	branch_block_stmt_2042/assign_stmt_2503_to_assign_stmt_2546/AND_u32_u32_2514_Sample/ra
      -- 
    ra_11746_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => AND_u32_u32_2514_inst_ack_0, ack => cp_elements(362)); -- 
    -- CP-element group 363 transition  input  output  bypass 
    -- predecessors 361 
    -- successors 365 
    -- members (10) 
      -- 	branch_block_stmt_2042/assign_stmt_2503_to_assign_stmt_2546/AND_u32_u32_2514_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2503_to_assign_stmt_2546/AND_u32_u32_2514_Update/$exit
      -- 	branch_block_stmt_2042/assign_stmt_2503_to_assign_stmt_2546/AND_u32_u32_2514_Update/ca
      -- 	branch_block_stmt_2042/assign_stmt_2503_to_assign_stmt_2546/ADD_u32_u32_2520_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_2503_to_assign_stmt_2546/R_iNsTr_141_2517_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_2503_to_assign_stmt_2546/R_iNsTr_141_2517_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2503_to_assign_stmt_2546/R_iNsTr_141_2517_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_2503_to_assign_stmt_2546/R_iNsTr_141_2517_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2503_to_assign_stmt_2546/ADD_u32_u32_2520_Sample/$entry
      -- 	branch_block_stmt_2042/assign_stmt_2503_to_assign_stmt_2546/ADD_u32_u32_2520_Sample/rr
      -- 
    ca_11751_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => AND_u32_u32_2514_inst_ack_1, ack => cp_elements(363)); -- 
    rr_11763_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(363), ack => ADD_u32_u32_2520_inst_req_0); -- 
    -- CP-element group 364 transition  output  bypass 
    -- predecessors 352 
    -- successors 366 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_2503_to_assign_stmt_2546/ADD_u32_u32_2520_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_2503_to_assign_stmt_2546/ADD_u32_u32_2520_Update/$entry
      -- 	branch_block_stmt_2042/assign_stmt_2503_to_assign_stmt_2546/ADD_u32_u32_2520_Update/cr
      -- 
    cp_elements(364) <= cp_elements(352);
    cr_11768_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(364), ack => ADD_u32_u32_2520_inst_req_1); -- 
    -- CP-element group 365 transition  input  bypass 
    -- predecessors 363 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_2503_to_assign_stmt_2546/ADD_u32_u32_2520_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2503_to_assign_stmt_2546/ADD_u32_u32_2520_Sample/$exit
      -- 	branch_block_stmt_2042/assign_stmt_2503_to_assign_stmt_2546/ADD_u32_u32_2520_Sample/ra
      -- 
    ra_11764_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u32_u32_2520_inst_ack_0, ack => cp_elements(365)); -- 
    -- CP-element group 366 transition  input  bypass 
    -- predecessors 364 
    -- successors 384 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_2503_to_assign_stmt_2546/ADD_u32_u32_2520_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2503_to_assign_stmt_2546/ADD_u32_u32_2520_Update/$exit
      -- 	branch_block_stmt_2042/assign_stmt_2503_to_assign_stmt_2546/ADD_u32_u32_2520_Update/ca
      -- 
    ca_11769_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u32_u32_2520_inst_ack_1, ack => cp_elements(366)); -- 
    -- CP-element group 367 transition  output  bypass 
    -- predecessors 352 
    -- successors 370 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_2503_to_assign_stmt_2546/AND_u32_u32_2526_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_2503_to_assign_stmt_2546/AND_u32_u32_2526_Update/$entry
      -- 	branch_block_stmt_2042/assign_stmt_2503_to_assign_stmt_2546/AND_u32_u32_2526_Update/cr
      -- 
    cp_elements(367) <= cp_elements(352);
    cr_11786_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(367), ack => AND_u32_u32_2526_inst_req_1); -- 
    -- CP-element group 368 transition  output  bypass 
    -- predecessors 352 
    -- successors 369 
    -- members (7) 
      -- 	branch_block_stmt_2042/assign_stmt_2503_to_assign_stmt_2546/AND_u32_u32_2526_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_2503_to_assign_stmt_2546/R_xx_xlcssa19_2523_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_2503_to_assign_stmt_2546/R_xx_xlcssa19_2523_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2503_to_assign_stmt_2546/R_xx_xlcssa19_2523_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_2503_to_assign_stmt_2546/R_xx_xlcssa19_2523_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2503_to_assign_stmt_2546/AND_u32_u32_2526_Sample/$entry
      -- 	branch_block_stmt_2042/assign_stmt_2503_to_assign_stmt_2546/AND_u32_u32_2526_Sample/rr
      -- 
    cp_elements(368) <= cp_elements(352);
    rr_11781_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(368), ack => AND_u32_u32_2526_inst_req_0); -- 
    -- CP-element group 369 transition  input  bypass 
    -- predecessors 368 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_2503_to_assign_stmt_2546/AND_u32_u32_2526_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2503_to_assign_stmt_2546/AND_u32_u32_2526_Sample/$exit
      -- 	branch_block_stmt_2042/assign_stmt_2503_to_assign_stmt_2546/AND_u32_u32_2526_Sample/ra
      -- 
    ra_11782_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => AND_u32_u32_2526_inst_ack_0, ack => cp_elements(369)); -- 
    -- CP-element group 370 transition  input  output  bypass 
    -- predecessors 367 
    -- successors 372 
    -- members (10) 
      -- 	branch_block_stmt_2042/assign_stmt_2503_to_assign_stmt_2546/AND_u32_u32_2526_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2503_to_assign_stmt_2546/AND_u32_u32_2526_Update/$exit
      -- 	branch_block_stmt_2042/assign_stmt_2503_to_assign_stmt_2546/AND_u32_u32_2526_Update/ca
      -- 	branch_block_stmt_2042/assign_stmt_2503_to_assign_stmt_2546/EQ_u32_u1_2532_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_2503_to_assign_stmt_2546/R_iNsTr_143_2529_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_2503_to_assign_stmt_2546/R_iNsTr_143_2529_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2503_to_assign_stmt_2546/R_iNsTr_143_2529_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_2503_to_assign_stmt_2546/R_iNsTr_143_2529_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2503_to_assign_stmt_2546/EQ_u32_u1_2532_Sample/$entry
      -- 	branch_block_stmt_2042/assign_stmt_2503_to_assign_stmt_2546/EQ_u32_u1_2532_Sample/rr
      -- 
    ca_11787_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => AND_u32_u32_2526_inst_ack_1, ack => cp_elements(370)); -- 
    rr_11799_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(370), ack => EQ_u32_u1_2532_inst_req_0); -- 
    -- CP-element group 371 transition  output  bypass 
    -- predecessors 352 
    -- successors 373 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_2503_to_assign_stmt_2546/EQ_u32_u1_2532_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_2503_to_assign_stmt_2546/EQ_u32_u1_2532_Update/$entry
      -- 	branch_block_stmt_2042/assign_stmt_2503_to_assign_stmt_2546/EQ_u32_u1_2532_Update/cr
      -- 
    cp_elements(371) <= cp_elements(352);
    cr_11804_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(371), ack => EQ_u32_u1_2532_inst_req_1); -- 
    -- CP-element group 372 transition  input  bypass 
    -- predecessors 370 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_2503_to_assign_stmt_2546/EQ_u32_u1_2532_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2503_to_assign_stmt_2546/EQ_u32_u1_2532_Sample/$exit
      -- 	branch_block_stmt_2042/assign_stmt_2503_to_assign_stmt_2546/EQ_u32_u1_2532_Sample/ra
      -- 
    ra_11800_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u32_u1_2532_inst_ack_0, ack => cp_elements(372)); -- 
    -- CP-element group 373 transition  input  bypass 
    -- predecessors 371 
    -- successors 380 
    -- members (7) 
      -- 	branch_block_stmt_2042/assign_stmt_2503_to_assign_stmt_2546/EQ_u32_u1_2532_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2503_to_assign_stmt_2546/EQ_u32_u1_2532_Update/$exit
      -- 	branch_block_stmt_2042/assign_stmt_2503_to_assign_stmt_2546/EQ_u32_u1_2532_Update/ca
      -- 	branch_block_stmt_2042/assign_stmt_2503_to_assign_stmt_2546/R_iNsTr_144_2543_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_2503_to_assign_stmt_2546/R_iNsTr_144_2543_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2503_to_assign_stmt_2546/R_iNsTr_144_2543_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_2503_to_assign_stmt_2546/R_iNsTr_144_2543_update_completed_
      -- 
    ca_11805_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u32_u1_2532_inst_ack_1, ack => cp_elements(373)); -- 
    -- CP-element group 374 transition  output  bypass 
    -- predecessors 352 
    -- successors 379 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_2503_to_assign_stmt_2546/NEQ_i32_u1_2540_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_2503_to_assign_stmt_2546/NEQ_i32_u1_2540_Update/$entry
      -- 	branch_block_stmt_2042/assign_stmt_2503_to_assign_stmt_2546/NEQ_i32_u1_2540_Update/cr
      -- 
    cp_elements(374) <= cp_elements(352);
    cr_11836_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(374), ack => NEQ_i32_u1_2540_inst_req_1); -- 
    -- CP-element group 375 transition  output  bypass 
    -- predecessors 352 
    -- successors 376 
    -- members (7) 
      -- 	branch_block_stmt_2042/assign_stmt_2503_to_assign_stmt_2546/type_cast_2536_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_2503_to_assign_stmt_2546/R_xx_xlcssa19_2535_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_2503_to_assign_stmt_2546/R_xx_xlcssa19_2535_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2503_to_assign_stmt_2546/R_xx_xlcssa19_2535_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_2503_to_assign_stmt_2546/R_xx_xlcssa19_2535_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2503_to_assign_stmt_2546/type_cast_2536_Sample/$entry
      -- 	branch_block_stmt_2042/assign_stmt_2503_to_assign_stmt_2546/type_cast_2536_Sample/rr
      -- 
    cp_elements(375) <= cp_elements(352);
    rr_11821_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(375), ack => type_cast_2536_inst_req_0); -- 
    -- CP-element group 376 transition  input  output  bypass 
    -- predecessors 375 
    -- successors 377 
    -- members (6) 
      -- 	branch_block_stmt_2042/assign_stmt_2503_to_assign_stmt_2546/type_cast_2536_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2503_to_assign_stmt_2546/type_cast_2536_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_2503_to_assign_stmt_2546/type_cast_2536_Sample/$exit
      -- 	branch_block_stmt_2042/assign_stmt_2503_to_assign_stmt_2546/type_cast_2536_Sample/ra
      -- 	branch_block_stmt_2042/assign_stmt_2503_to_assign_stmt_2546/type_cast_2536_Update/$entry
      -- 	branch_block_stmt_2042/assign_stmt_2503_to_assign_stmt_2546/type_cast_2536_Update/cr
      -- 
    ra_11822_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2536_inst_ack_0, ack => cp_elements(376)); -- 
    cr_11826_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(376), ack => type_cast_2536_inst_req_1); -- 
    -- CP-element group 377 transition  input  output  bypass 
    -- predecessors 376 
    -- successors 378 
    -- members (6) 
      -- 	branch_block_stmt_2042/assign_stmt_2503_to_assign_stmt_2546/NEQ_i32_u1_2540_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_2503_to_assign_stmt_2546/type_cast_2536_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2503_to_assign_stmt_2546/type_cast_2536_Update/$exit
      -- 	branch_block_stmt_2042/assign_stmt_2503_to_assign_stmt_2546/type_cast_2536_Update/ca
      -- 	branch_block_stmt_2042/assign_stmt_2503_to_assign_stmt_2546/NEQ_i32_u1_2540_Sample/$entry
      -- 	branch_block_stmt_2042/assign_stmt_2503_to_assign_stmt_2546/NEQ_i32_u1_2540_Sample/rr
      -- 
    ca_11827_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2536_inst_ack_1, ack => cp_elements(377)); -- 
    rr_11831_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(377), ack => NEQ_i32_u1_2540_inst_req_0); -- 
    -- CP-element group 378 transition  input  bypass 
    -- predecessors 377 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_2503_to_assign_stmt_2546/NEQ_i32_u1_2540_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2503_to_assign_stmt_2546/NEQ_i32_u1_2540_Sample/$exit
      -- 	branch_block_stmt_2042/assign_stmt_2503_to_assign_stmt_2546/NEQ_i32_u1_2540_Sample/ra
      -- 
    ra_11832_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => NEQ_i32_u1_2540_inst_ack_0, ack => cp_elements(378)); -- 
    -- CP-element group 379 transition  input  bypass 
    -- predecessors 374 
    -- successors 380 
    -- members (7) 
      -- 	branch_block_stmt_2042/assign_stmt_2503_to_assign_stmt_2546/NEQ_i32_u1_2540_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2503_to_assign_stmt_2546/NEQ_i32_u1_2540_Update/$exit
      -- 	branch_block_stmt_2042/assign_stmt_2503_to_assign_stmt_2546/NEQ_i32_u1_2540_Update/ca
      -- 	branch_block_stmt_2042/assign_stmt_2503_to_assign_stmt_2546/R_iNsTr_145_2544_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_2503_to_assign_stmt_2546/R_iNsTr_145_2544_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2503_to_assign_stmt_2546/R_iNsTr_145_2544_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_2503_to_assign_stmt_2546/R_iNsTr_145_2544_update_completed_
      -- 
    ca_11837_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => NEQ_i32_u1_2540_inst_ack_1, ack => cp_elements(379)); -- 
    -- CP-element group 380 join  transition  output  bypass 
    -- predecessors 373 379 
    -- successors 382 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_2503_to_assign_stmt_2546/AND_u1_u1_2545_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_2503_to_assign_stmt_2546/AND_u1_u1_2545_Sample/$entry
      -- 	branch_block_stmt_2042/assign_stmt_2503_to_assign_stmt_2546/AND_u1_u1_2545_Sample/rr
      -- 
    cp_element_group_380: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 20) := "cp_element_group_380"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(373) & cp_elements(379);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(380), clk => clk, reset => reset); --
    end block;
    rr_11853_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(380), ack => AND_u1_u1_2545_inst_req_0); -- 
    -- CP-element group 381 transition  output  bypass 
    -- predecessors 352 
    -- successors 383 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_2503_to_assign_stmt_2546/AND_u1_u1_2545_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_2503_to_assign_stmt_2546/AND_u1_u1_2545_Update/$entry
      -- 	branch_block_stmt_2042/assign_stmt_2503_to_assign_stmt_2546/AND_u1_u1_2545_Update/cr
      -- 
    cp_elements(381) <= cp_elements(352);
    cr_11858_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(381), ack => AND_u1_u1_2545_inst_req_1); -- 
    -- CP-element group 382 transition  input  bypass 
    -- predecessors 380 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_2503_to_assign_stmt_2546/AND_u1_u1_2545_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2503_to_assign_stmt_2546/AND_u1_u1_2545_Sample/$exit
      -- 	branch_block_stmt_2042/assign_stmt_2503_to_assign_stmt_2546/AND_u1_u1_2545_Sample/ra
      -- 
    ra_11854_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => AND_u1_u1_2545_inst_ack_0, ack => cp_elements(382)); -- 
    -- CP-element group 383 transition  input  bypass 
    -- predecessors 381 
    -- successors 384 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_2503_to_assign_stmt_2546/AND_u1_u1_2545_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2503_to_assign_stmt_2546/AND_u1_u1_2545_Update/$exit
      -- 	branch_block_stmt_2042/assign_stmt_2503_to_assign_stmt_2546/AND_u1_u1_2545_Update/ca
      -- 
    ca_11859_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => AND_u1_u1_2545_inst_ack_1, ack => cp_elements(383)); -- 
    -- CP-element group 384 join  transition  bypass 
    -- predecessors 360 366 383 
    -- successors 20 
    -- members (1) 
      -- 	branch_block_stmt_2042/assign_stmt_2503_to_assign_stmt_2546/$exit
      -- 
    cp_element_group_384: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 20) := "cp_element_group_384"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= cp_elements(360) & cp_elements(366) & cp_elements(383);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(384), clk => clk, reset => reset); --
    end block;
    -- CP-element group 385 transition  place  dead  bypass 
    -- predecessors 20 
    -- successors 21 
    -- members (8) 
      -- 	branch_block_stmt_2042/if_stmt_2547__exit__
      -- 	branch_block_stmt_2042/merge_stmt_2553__entry__
      -- 	branch_block_stmt_2042/if_stmt_2547_dead_link/$entry
      -- 	branch_block_stmt_2042/if_stmt_2547_dead_link/$exit
      -- 	branch_block_stmt_2042/if_stmt_2547_dead_link/dead_transition
      -- 	branch_block_stmt_2042/merge_stmt_2553_dead_link/$entry
      -- 	branch_block_stmt_2042/merge_stmt_2553_dead_link/$exit
      -- 	branch_block_stmt_2042/merge_stmt_2553_dead_link/dead_transition
      -- 
    cp_elements(385) <= false;
    -- CP-element group 386 transition  output  bypass 
    -- predecessors 20 
    -- successors 387 
    -- members (3) 
      -- 	branch_block_stmt_2042/if_stmt_2547_eval_test/$entry
      -- 	branch_block_stmt_2042/if_stmt_2547_eval_test/$exit
      -- 	branch_block_stmt_2042/if_stmt_2547_eval_test/branch_req
      -- 
    cp_elements(386) <= cp_elements(20);
    branch_req_11867_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(386), ack => if_stmt_2547_branch_req_0); -- 
    -- CP-element group 387 branch  place  bypass 
    -- predecessors 386 
    -- successors 388 390 
    -- members (1) 
      -- 	branch_block_stmt_2042/R_orx_xcond11x_xix_xi40_2548_place
      -- 
    cp_elements(387) <= cp_elements(386);
    -- CP-element group 388 transition  bypass 
    -- predecessors 387 
    -- successors 389 
    -- members (1) 
      -- 	branch_block_stmt_2042/if_stmt_2547_if_link/$entry
      -- 
    cp_elements(388) <= cp_elements(387);
    -- CP-element group 389 transition  place  input  bypass 
    -- predecessors 388 
    -- successors 21 
    -- members (9) 
      -- 	branch_block_stmt_2042/if_stmt_2547_if_link/$exit
      -- 	branch_block_stmt_2042/if_stmt_2547_if_link/if_choice_transition
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xpreheaderx_xix_xi41_udiv32x_xexitx_xix_xi45x_xpreheader
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xpreheaderx_xix_xi41_udiv32x_xexitx_xix_xi45x_xpreheader_PhiReq/$entry
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xpreheaderx_xix_xi41_udiv32x_xexitx_xix_xi45x_xpreheader_PhiReq/$exit
      -- 	branch_block_stmt_2042/merge_stmt_2553_PhiReqMerge
      -- 	branch_block_stmt_2042/merge_stmt_2553_PhiAck/$entry
      -- 	branch_block_stmt_2042/merge_stmt_2553_PhiAck/$exit
      -- 	branch_block_stmt_2042/merge_stmt_2553_PhiAck/dummy
      -- 
    if_choice_transition_11872_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2547_branch_ack_1, ack => cp_elements(389)); -- 
    -- CP-element group 390 transition  bypass 
    -- predecessors 387 
    -- successors 391 
    -- members (1) 
      -- 	branch_block_stmt_2042/if_stmt_2547_else_link/$entry
      -- 
    cp_elements(390) <= cp_elements(387);
    -- CP-element group 391 transition  place  input  bypass 
    -- predecessors 390 
    -- successors 1594 
    -- members (3) 
      -- 	branch_block_stmt_2042/if_stmt_2547_else_link/$exit
      -- 	branch_block_stmt_2042/if_stmt_2547_else_link/else_choice_transition
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xpreheaderx_xix_xi41_xx_xcritedgex_xix_xi52
      -- 
    else_choice_transition_11876_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2547_branch_ack_0, ack => cp_elements(391)); -- 
    -- CP-element group 392 fork  transition  bypass 
    -- predecessors 22 
    -- successors 393 394 397 401 404 411 414 415 
    -- members (1) 
      -- 	branch_block_stmt_2042/assign_stmt_2575_to_assign_stmt_2606/$entry
      -- 
    cp_elements(392) <= cp_elements(22);
    -- CP-element group 393 transition  output  bypass 
    -- predecessors 392 
    -- successors 396 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_2575_to_assign_stmt_2606/SHL_u32_u32_2574_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_2575_to_assign_stmt_2606/SHL_u32_u32_2574_Update/$entry
      -- 	branch_block_stmt_2042/assign_stmt_2575_to_assign_stmt_2606/SHL_u32_u32_2574_Update/cr
      -- 
    cp_elements(393) <= cp_elements(392);
    cr_11898_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(393), ack => SHL_u32_u32_2574_inst_req_1); -- 
    -- CP-element group 394 transition  output  bypass 
    -- predecessors 392 
    -- successors 395 
    -- members (7) 
      -- 	branch_block_stmt_2042/assign_stmt_2575_to_assign_stmt_2606/SHL_u32_u32_2574_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_2575_to_assign_stmt_2606/R_tempx_x012x_xix_xi42_2571_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_2575_to_assign_stmt_2606/R_tempx_x012x_xix_xi42_2571_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2575_to_assign_stmt_2606/R_tempx_x012x_xix_xi42_2571_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_2575_to_assign_stmt_2606/R_tempx_x012x_xix_xi42_2571_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2575_to_assign_stmt_2606/SHL_u32_u32_2574_Sample/$entry
      -- 	branch_block_stmt_2042/assign_stmt_2575_to_assign_stmt_2606/SHL_u32_u32_2574_Sample/rr
      -- 
    cp_elements(394) <= cp_elements(392);
    rr_11893_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(394), ack => SHL_u32_u32_2574_inst_req_0); -- 
    -- CP-element group 395 transition  input  bypass 
    -- predecessors 394 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_2575_to_assign_stmt_2606/SHL_u32_u32_2574_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2575_to_assign_stmt_2606/SHL_u32_u32_2574_Sample/$exit
      -- 	branch_block_stmt_2042/assign_stmt_2575_to_assign_stmt_2606/SHL_u32_u32_2574_Sample/ra
      -- 
    ra_11894_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => SHL_u32_u32_2574_inst_ack_0, ack => cp_elements(395)); -- 
    -- CP-element group 396 fork  transition  input  bypass 
    -- predecessors 393 
    -- successors 398 405 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_2575_to_assign_stmt_2606/SHL_u32_u32_2574_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2575_to_assign_stmt_2606/SHL_u32_u32_2574_Update/$exit
      -- 	branch_block_stmt_2042/assign_stmt_2575_to_assign_stmt_2606/SHL_u32_u32_2574_Update/ca
      -- 
    ca_11899_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => SHL_u32_u32_2574_inst_ack_1, ack => cp_elements(396)); -- 
    -- CP-element group 397 transition  output  bypass 
    -- predecessors 392 
    -- successors 400 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_2575_to_assign_stmt_2606/AND_u32_u32_2580_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_2575_to_assign_stmt_2606/AND_u32_u32_2580_Update/$entry
      -- 	branch_block_stmt_2042/assign_stmt_2575_to_assign_stmt_2606/AND_u32_u32_2580_Update/cr
      -- 
    cp_elements(397) <= cp_elements(392);
    cr_11916_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(397), ack => AND_u32_u32_2580_inst_req_1); -- 
    -- CP-element group 398 transition  output  bypass 
    -- predecessors 396 
    -- successors 399 
    -- members (7) 
      -- 	branch_block_stmt_2042/assign_stmt_2575_to_assign_stmt_2606/AND_u32_u32_2580_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_2575_to_assign_stmt_2606/R_iNsTr_206_2577_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_2575_to_assign_stmt_2606/R_iNsTr_206_2577_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2575_to_assign_stmt_2606/R_iNsTr_206_2577_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_2575_to_assign_stmt_2606/R_iNsTr_206_2577_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2575_to_assign_stmt_2606/AND_u32_u32_2580_Sample/$entry
      -- 	branch_block_stmt_2042/assign_stmt_2575_to_assign_stmt_2606/AND_u32_u32_2580_Sample/rr
      -- 
    cp_elements(398) <= cp_elements(396);
    rr_11911_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(398), ack => AND_u32_u32_2580_inst_req_0); -- 
    -- CP-element group 399 transition  input  bypass 
    -- predecessors 398 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_2575_to_assign_stmt_2606/AND_u32_u32_2580_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2575_to_assign_stmt_2606/AND_u32_u32_2580_Sample/$exit
      -- 	branch_block_stmt_2042/assign_stmt_2575_to_assign_stmt_2606/AND_u32_u32_2580_Sample/ra
      -- 
    ra_11912_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => AND_u32_u32_2580_inst_ack_0, ack => cp_elements(399)); -- 
    -- CP-element group 400 transition  input  output  bypass 
    -- predecessors 397 
    -- successors 402 
    -- members (10) 
      -- 	branch_block_stmt_2042/assign_stmt_2575_to_assign_stmt_2606/AND_u32_u32_2580_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2575_to_assign_stmt_2606/AND_u32_u32_2580_Update/$exit
      -- 	branch_block_stmt_2042/assign_stmt_2575_to_assign_stmt_2606/AND_u32_u32_2580_Update/ca
      -- 	branch_block_stmt_2042/assign_stmt_2575_to_assign_stmt_2606/EQ_u32_u1_2586_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_2575_to_assign_stmt_2606/R_iNsTr_207_2583_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_2575_to_assign_stmt_2606/R_iNsTr_207_2583_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2575_to_assign_stmt_2606/R_iNsTr_207_2583_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_2575_to_assign_stmt_2606/R_iNsTr_207_2583_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2575_to_assign_stmt_2606/EQ_u32_u1_2586_Sample/$entry
      -- 	branch_block_stmt_2042/assign_stmt_2575_to_assign_stmt_2606/EQ_u32_u1_2586_Sample/rr
      -- 
    ca_11917_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => AND_u32_u32_2580_inst_ack_1, ack => cp_elements(400)); -- 
    rr_11929_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(400), ack => EQ_u32_u1_2586_inst_req_0); -- 
    -- CP-element group 401 transition  output  bypass 
    -- predecessors 392 
    -- successors 403 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_2575_to_assign_stmt_2606/EQ_u32_u1_2586_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_2575_to_assign_stmt_2606/EQ_u32_u1_2586_Update/$entry
      -- 	branch_block_stmt_2042/assign_stmt_2575_to_assign_stmt_2606/EQ_u32_u1_2586_Update/cr
      -- 
    cp_elements(401) <= cp_elements(392);
    cr_11934_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(401), ack => EQ_u32_u1_2586_inst_req_1); -- 
    -- CP-element group 402 transition  input  bypass 
    -- predecessors 400 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_2575_to_assign_stmt_2606/EQ_u32_u1_2586_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2575_to_assign_stmt_2606/EQ_u32_u1_2586_Sample/$exit
      -- 	branch_block_stmt_2042/assign_stmt_2575_to_assign_stmt_2606/EQ_u32_u1_2586_Sample/ra
      -- 
    ra_11930_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u32_u1_2586_inst_ack_0, ack => cp_elements(402)); -- 
    -- CP-element group 403 transition  input  bypass 
    -- predecessors 401 
    -- successors 410 
    -- members (7) 
      -- 	branch_block_stmt_2042/assign_stmt_2575_to_assign_stmt_2606/EQ_u32_u1_2586_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2575_to_assign_stmt_2606/EQ_u32_u1_2586_Update/$exit
      -- 	branch_block_stmt_2042/assign_stmt_2575_to_assign_stmt_2606/EQ_u32_u1_2586_Update/ca
      -- 	branch_block_stmt_2042/assign_stmt_2575_to_assign_stmt_2606/R_iNsTr_208_2597_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_2575_to_assign_stmt_2606/R_iNsTr_208_2597_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2575_to_assign_stmt_2606/R_iNsTr_208_2597_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_2575_to_assign_stmt_2606/R_iNsTr_208_2597_update_completed_
      -- 
    ca_11935_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u32_u1_2586_inst_ack_1, ack => cp_elements(403)); -- 
    -- CP-element group 404 transition  output  bypass 
    -- predecessors 392 
    -- successors 409 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_2575_to_assign_stmt_2606/NEQ_i32_u1_2594_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_2575_to_assign_stmt_2606/NEQ_i32_u1_2594_Update/$entry
      -- 	branch_block_stmt_2042/assign_stmt_2575_to_assign_stmt_2606/NEQ_i32_u1_2594_Update/cr
      -- 
    cp_elements(404) <= cp_elements(392);
    cr_11966_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(404), ack => NEQ_i32_u1_2594_inst_req_1); -- 
    -- CP-element group 405 transition  output  bypass 
    -- predecessors 396 
    -- successors 406 
    -- members (7) 
      -- 	branch_block_stmt_2042/assign_stmt_2575_to_assign_stmt_2606/type_cast_2590_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_2575_to_assign_stmt_2606/R_iNsTr_206_2589_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_2575_to_assign_stmt_2606/R_iNsTr_206_2589_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2575_to_assign_stmt_2606/R_iNsTr_206_2589_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_2575_to_assign_stmt_2606/R_iNsTr_206_2589_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2575_to_assign_stmt_2606/type_cast_2590_Sample/$entry
      -- 	branch_block_stmt_2042/assign_stmt_2575_to_assign_stmt_2606/type_cast_2590_Sample/rr
      -- 
    cp_elements(405) <= cp_elements(396);
    rr_11951_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(405), ack => type_cast_2590_inst_req_0); -- 
    -- CP-element group 406 transition  input  output  bypass 
    -- predecessors 405 
    -- successors 407 
    -- members (6) 
      -- 	branch_block_stmt_2042/assign_stmt_2575_to_assign_stmt_2606/type_cast_2590_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2575_to_assign_stmt_2606/type_cast_2590_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_2575_to_assign_stmt_2606/type_cast_2590_Sample/$exit
      -- 	branch_block_stmt_2042/assign_stmt_2575_to_assign_stmt_2606/type_cast_2590_Sample/ra
      -- 	branch_block_stmt_2042/assign_stmt_2575_to_assign_stmt_2606/type_cast_2590_Update/$entry
      -- 	branch_block_stmt_2042/assign_stmt_2575_to_assign_stmt_2606/type_cast_2590_Update/cr
      -- 
    ra_11952_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2590_inst_ack_0, ack => cp_elements(406)); -- 
    cr_11956_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(406), ack => type_cast_2590_inst_req_1); -- 
    -- CP-element group 407 transition  input  output  bypass 
    -- predecessors 406 
    -- successors 408 
    -- members (6) 
      -- 	branch_block_stmt_2042/assign_stmt_2575_to_assign_stmt_2606/NEQ_i32_u1_2594_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_2575_to_assign_stmt_2606/type_cast_2590_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2575_to_assign_stmt_2606/type_cast_2590_Update/$exit
      -- 	branch_block_stmt_2042/assign_stmt_2575_to_assign_stmt_2606/type_cast_2590_Update/ca
      -- 	branch_block_stmt_2042/assign_stmt_2575_to_assign_stmt_2606/NEQ_i32_u1_2594_Sample/$entry
      -- 	branch_block_stmt_2042/assign_stmt_2575_to_assign_stmt_2606/NEQ_i32_u1_2594_Sample/rr
      -- 
    ca_11957_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2590_inst_ack_1, ack => cp_elements(407)); -- 
    rr_11961_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(407), ack => NEQ_i32_u1_2594_inst_req_0); -- 
    -- CP-element group 408 transition  input  bypass 
    -- predecessors 407 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_2575_to_assign_stmt_2606/NEQ_i32_u1_2594_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2575_to_assign_stmt_2606/NEQ_i32_u1_2594_Sample/$exit
      -- 	branch_block_stmt_2042/assign_stmt_2575_to_assign_stmt_2606/NEQ_i32_u1_2594_Sample/ra
      -- 
    ra_11962_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => NEQ_i32_u1_2594_inst_ack_0, ack => cp_elements(408)); -- 
    -- CP-element group 409 transition  input  bypass 
    -- predecessors 404 
    -- successors 410 
    -- members (7) 
      -- 	branch_block_stmt_2042/assign_stmt_2575_to_assign_stmt_2606/NEQ_i32_u1_2594_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2575_to_assign_stmt_2606/NEQ_i32_u1_2594_Update/$exit
      -- 	branch_block_stmt_2042/assign_stmt_2575_to_assign_stmt_2606/NEQ_i32_u1_2594_Update/ca
      -- 	branch_block_stmt_2042/assign_stmt_2575_to_assign_stmt_2606/R_iNsTr_209_2598_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_2575_to_assign_stmt_2606/R_iNsTr_209_2598_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2575_to_assign_stmt_2606/R_iNsTr_209_2598_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_2575_to_assign_stmt_2606/R_iNsTr_209_2598_update_completed_
      -- 
    ca_11967_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => NEQ_i32_u1_2594_inst_ack_1, ack => cp_elements(409)); -- 
    -- CP-element group 410 join  transition  output  bypass 
    -- predecessors 403 409 
    -- successors 412 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_2575_to_assign_stmt_2606/AND_u1_u1_2599_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_2575_to_assign_stmt_2606/AND_u1_u1_2599_Sample/$entry
      -- 	branch_block_stmt_2042/assign_stmt_2575_to_assign_stmt_2606/AND_u1_u1_2599_Sample/rr
      -- 
    cp_element_group_410: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 20) := "cp_element_group_410"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(403) & cp_elements(409);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(410), clk => clk, reset => reset); --
    end block;
    rr_11983_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(410), ack => AND_u1_u1_2599_inst_req_0); -- 
    -- CP-element group 411 transition  output  bypass 
    -- predecessors 392 
    -- successors 413 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_2575_to_assign_stmt_2606/AND_u1_u1_2599_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_2575_to_assign_stmt_2606/AND_u1_u1_2599_Update/$entry
      -- 	branch_block_stmt_2042/assign_stmt_2575_to_assign_stmt_2606/AND_u1_u1_2599_Update/cr
      -- 
    cp_elements(411) <= cp_elements(392);
    cr_11988_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(411), ack => AND_u1_u1_2599_inst_req_1); -- 
    -- CP-element group 412 transition  input  bypass 
    -- predecessors 410 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_2575_to_assign_stmt_2606/AND_u1_u1_2599_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2575_to_assign_stmt_2606/AND_u1_u1_2599_Sample/$exit
      -- 	branch_block_stmt_2042/assign_stmt_2575_to_assign_stmt_2606/AND_u1_u1_2599_Sample/ra
      -- 
    ra_11984_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => AND_u1_u1_2599_inst_ack_0, ack => cp_elements(412)); -- 
    -- CP-element group 413 transition  input  bypass 
    -- predecessors 411 
    -- successors 418 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_2575_to_assign_stmt_2606/AND_u1_u1_2599_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2575_to_assign_stmt_2606/AND_u1_u1_2599_Update/$exit
      -- 	branch_block_stmt_2042/assign_stmt_2575_to_assign_stmt_2606/AND_u1_u1_2599_Update/ca
      -- 
    ca_11989_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => AND_u1_u1_2599_inst_ack_1, ack => cp_elements(413)); -- 
    -- CP-element group 414 transition  output  bypass 
    -- predecessors 392 
    -- successors 417 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_2575_to_assign_stmt_2606/ADD_u32_u32_2605_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_2575_to_assign_stmt_2606/ADD_u32_u32_2605_Update/$entry
      -- 	branch_block_stmt_2042/assign_stmt_2575_to_assign_stmt_2606/ADD_u32_u32_2605_Update/cr
      -- 
    cp_elements(414) <= cp_elements(392);
    cr_12006_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(414), ack => ADD_u32_u32_2605_inst_req_1); -- 
    -- CP-element group 415 transition  output  bypass 
    -- predecessors 392 
    -- successors 416 
    -- members (7) 
      -- 	branch_block_stmt_2042/assign_stmt_2575_to_assign_stmt_2606/ADD_u32_u32_2605_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_2575_to_assign_stmt_2606/R_iNsTr_205_2602_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_2575_to_assign_stmt_2606/R_iNsTr_205_2602_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2575_to_assign_stmt_2606/R_iNsTr_205_2602_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_2575_to_assign_stmt_2606/R_iNsTr_205_2602_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2575_to_assign_stmt_2606/ADD_u32_u32_2605_Sample/$entry
      -- 	branch_block_stmt_2042/assign_stmt_2575_to_assign_stmt_2606/ADD_u32_u32_2605_Sample/rr
      -- 
    cp_elements(415) <= cp_elements(392);
    rr_12001_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(415), ack => ADD_u32_u32_2605_inst_req_0); -- 
    -- CP-element group 416 transition  input  bypass 
    -- predecessors 415 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_2575_to_assign_stmt_2606/ADD_u32_u32_2605_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2575_to_assign_stmt_2606/ADD_u32_u32_2605_Sample/$exit
      -- 	branch_block_stmt_2042/assign_stmt_2575_to_assign_stmt_2606/ADD_u32_u32_2605_Sample/ra
      -- 
    ra_12002_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u32_u32_2605_inst_ack_0, ack => cp_elements(416)); -- 
    -- CP-element group 417 transition  input  bypass 
    -- predecessors 414 
    -- successors 418 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_2575_to_assign_stmt_2606/ADD_u32_u32_2605_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2575_to_assign_stmt_2606/ADD_u32_u32_2605_Update/$exit
      -- 	branch_block_stmt_2042/assign_stmt_2575_to_assign_stmt_2606/ADD_u32_u32_2605_Update/ca
      -- 
    ca_12007_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u32_u32_2605_inst_ack_1, ack => cp_elements(417)); -- 
    -- CP-element group 418 join  transition  bypass 
    -- predecessors 413 417 
    -- successors 23 
    -- members (1) 
      -- 	branch_block_stmt_2042/assign_stmt_2575_to_assign_stmt_2606/$exit
      -- 
    cp_element_group_418: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 20) := "cp_element_group_418"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(413) & cp_elements(417);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(418), clk => clk, reset => reset); --
    end block;
    -- CP-element group 419 transition  place  dead  bypass 
    -- predecessors 23 
    -- successors 24 
    -- members (8) 
      -- 	branch_block_stmt_2042/if_stmt_2607__exit__
      -- 	branch_block_stmt_2042/merge_stmt_2613__entry__
      -- 	branch_block_stmt_2042/if_stmt_2607_dead_link/$entry
      -- 	branch_block_stmt_2042/if_stmt_2607_dead_link/$exit
      -- 	branch_block_stmt_2042/if_stmt_2607_dead_link/dead_transition
      -- 	branch_block_stmt_2042/merge_stmt_2613_dead_link/$entry
      -- 	branch_block_stmt_2042/merge_stmt_2613_dead_link/$exit
      -- 	branch_block_stmt_2042/merge_stmt_2613_dead_link/dead_transition
      -- 
    cp_elements(419) <= false;
    -- CP-element group 420 transition  output  bypass 
    -- predecessors 23 
    -- successors 421 
    -- members (3) 
      -- 	branch_block_stmt_2042/if_stmt_2607_eval_test/$entry
      -- 	branch_block_stmt_2042/if_stmt_2607_eval_test/$exit
      -- 	branch_block_stmt_2042/if_stmt_2607_eval_test/branch_req
      -- 
    cp_elements(420) <= cp_elements(23);
    branch_req_12015_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(420), ack => if_stmt_2607_branch_req_0); -- 
    -- CP-element group 421 branch  place  bypass 
    -- predecessors 420 
    -- successors 422 424 
    -- members (1) 
      -- 	branch_block_stmt_2042/R_orx_xcondx_xix_xi43_2608_place
      -- 
    cp_elements(421) <= cp_elements(420);
    -- CP-element group 422 transition  bypass 
    -- predecessors 421 
    -- successors 423 
    -- members (1) 
      -- 	branch_block_stmt_2042/if_stmt_2607_if_link/$entry
      -- 
    cp_elements(422) <= cp_elements(421);
    -- CP-element group 423 transition  place  input  bypass 
    -- predecessors 422 
    -- successors 1532 
    -- members (3) 
      -- 	branch_block_stmt_2042/if_stmt_2607_if_link/$exit
      -- 	branch_block_stmt_2042/if_stmt_2607_if_link/if_choice_transition
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi45_udiv32x_xexitx_xix_xi45
      -- 
    if_choice_transition_12020_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2607_branch_ack_1, ack => cp_elements(423)); -- 
    -- CP-element group 424 transition  bypass 
    -- predecessors 421 
    -- successors 425 
    -- members (1) 
      -- 	branch_block_stmt_2042/if_stmt_2607_else_link/$entry
      -- 
    cp_elements(424) <= cp_elements(421);
    -- CP-element group 425 transition  place  input  bypass 
    -- predecessors 424 
    -- successors 1575 
    -- members (3) 
      -- 	branch_block_stmt_2042/if_stmt_2607_else_link/$exit
      -- 	branch_block_stmt_2042/if_stmt_2607_else_link/else_choice_transition
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi45_udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi48
      -- 
    else_choice_transition_12024_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2607_branch_ack_0, ack => cp_elements(425)); -- 
    -- CP-element group 426 fork  transition  bypass 
    -- predecessors 24 
    -- successors 427 428 432 433 
    -- members (1) 
      -- 	branch_block_stmt_2042/assign_stmt_2628_to_assign_stmt_2633/$entry
      -- 
    cp_elements(426) <= cp_elements(24);
    -- CP-element group 427 transition  output  bypass 
    -- predecessors 426 
    -- successors 430 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_2628_to_assign_stmt_2633/ADD_u32_u32_2627_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_2628_to_assign_stmt_2633/ADD_u32_u32_2627_Update/$entry
      -- 	branch_block_stmt_2042/assign_stmt_2628_to_assign_stmt_2633/ADD_u32_u32_2627_Update/cr
      -- 
    cp_elements(427) <= cp_elements(426);
    cr_12046_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(427), ack => ADD_u32_u32_2627_inst_req_1); -- 
    -- CP-element group 428 transition  output  bypass 
    -- predecessors 426 
    -- successors 429 
    -- members (7) 
      -- 	branch_block_stmt_2042/assign_stmt_2628_to_assign_stmt_2633/ADD_u32_u32_2627_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_2628_to_assign_stmt_2633/R_iNsTr_141_2624_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_2628_to_assign_stmt_2633/R_iNsTr_141_2624_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2628_to_assign_stmt_2633/R_iNsTr_141_2624_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_2628_to_assign_stmt_2633/R_iNsTr_141_2624_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2628_to_assign_stmt_2633/ADD_u32_u32_2627_Sample/$entry
      -- 	branch_block_stmt_2042/assign_stmt_2628_to_assign_stmt_2633/ADD_u32_u32_2627_Sample/rr
      -- 
    cp_elements(428) <= cp_elements(426);
    rr_12041_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(428), ack => ADD_u32_u32_2627_inst_req_0); -- 
    -- CP-element group 429 transition  input  bypass 
    -- predecessors 428 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_2628_to_assign_stmt_2633/ADD_u32_u32_2627_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2628_to_assign_stmt_2633/ADD_u32_u32_2627_Sample/$exit
      -- 	branch_block_stmt_2042/assign_stmt_2628_to_assign_stmt_2633/ADD_u32_u32_2627_Sample/ra
      -- 
    ra_12042_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u32_u32_2627_inst_ack_0, ack => cp_elements(429)); -- 
    -- CP-element group 430 transition  input  bypass 
    -- predecessors 427 
    -- successors 431 
    -- members (7) 
      -- 	branch_block_stmt_2042/assign_stmt_2628_to_assign_stmt_2633/ADD_u32_u32_2627_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2628_to_assign_stmt_2633/ADD_u32_u32_2627_Update/$exit
      -- 	branch_block_stmt_2042/assign_stmt_2628_to_assign_stmt_2633/ADD_u32_u32_2627_Update/ca
      -- 	branch_block_stmt_2042/assign_stmt_2628_to_assign_stmt_2633/R_tmp25x_xix_xi46_2630_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_2628_to_assign_stmt_2633/R_tmp25x_xix_xi46_2630_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2628_to_assign_stmt_2633/R_tmp25x_xix_xi46_2630_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_2628_to_assign_stmt_2633/R_tmp25x_xix_xi46_2630_update_completed_
      -- 
    ca_12047_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u32_u32_2627_inst_ack_1, ack => cp_elements(430)); -- 
    -- CP-element group 431 join  transition  output  bypass 
    -- predecessors 430 433 
    -- successors 434 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_2628_to_assign_stmt_2633/SUB_u32_u32_2632_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_2628_to_assign_stmt_2633/SUB_u32_u32_2632_Sample/$entry
      -- 	branch_block_stmt_2042/assign_stmt_2628_to_assign_stmt_2633/SUB_u32_u32_2632_Sample/rr
      -- 
    cp_element_group_431: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 20) := "cp_element_group_431"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(430) & cp_elements(433);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(431), clk => clk, reset => reset); --
    end block;
    rr_12063_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(431), ack => SUB_u32_u32_2632_inst_req_0); -- 
    -- CP-element group 432 transition  output  bypass 
    -- predecessors 426 
    -- successors 435 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_2628_to_assign_stmt_2633/SUB_u32_u32_2632_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_2628_to_assign_stmt_2633/SUB_u32_u32_2632_Update/$entry
      -- 	branch_block_stmt_2042/assign_stmt_2628_to_assign_stmt_2633/SUB_u32_u32_2632_Update/cr
      -- 
    cp_elements(432) <= cp_elements(426);
    cr_12068_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(432), ack => SUB_u32_u32_2632_inst_req_1); -- 
    -- CP-element group 433 transition  bypass 
    -- predecessors 426 
    -- successors 431 
    -- members (4) 
      -- 	branch_block_stmt_2042/assign_stmt_2628_to_assign_stmt_2633/R_xx_xlcssa15_2631_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_2628_to_assign_stmt_2633/R_xx_xlcssa15_2631_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2628_to_assign_stmt_2633/R_xx_xlcssa15_2631_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_2628_to_assign_stmt_2633/R_xx_xlcssa15_2631_update_completed_
      -- 
    cp_elements(433) <= cp_elements(426);
    -- CP-element group 434 transition  input  bypass 
    -- predecessors 431 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_2628_to_assign_stmt_2633/SUB_u32_u32_2632_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2628_to_assign_stmt_2633/SUB_u32_u32_2632_Sample/$exit
      -- 	branch_block_stmt_2042/assign_stmt_2628_to_assign_stmt_2633/SUB_u32_u32_2632_Sample/ra
      -- 
    ra_12064_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => SUB_u32_u32_2632_inst_ack_0, ack => cp_elements(434)); -- 
    -- CP-element group 435 transition  place  input  bypass 
    -- predecessors 432 
    -- successors 1620 
    -- members (6) 
      -- 	branch_block_stmt_2042/assign_stmt_2628_to_assign_stmt_2633__exit__
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi48_xx_xcritedgex_xix_xi52
      -- 	branch_block_stmt_2042/assign_stmt_2628_to_assign_stmt_2633/$exit
      -- 	branch_block_stmt_2042/assign_stmt_2628_to_assign_stmt_2633/SUB_u32_u32_2632_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2628_to_assign_stmt_2633/SUB_u32_u32_2632_Update/$exit
      -- 	branch_block_stmt_2042/assign_stmt_2628_to_assign_stmt_2633/SUB_u32_u32_2632_Update/ca
      -- 
    ca_12069_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => SUB_u32_u32_2632_inst_ack_1, ack => cp_elements(435)); -- 
    -- CP-element group 436 fork  transition  bypass 
    -- predecessors 25 
    -- successors 437 438 441 442 445 449 450 454 457 
    -- members (1) 
      -- 	branch_block_stmt_2042/assign_stmt_2654_to_assign_stmt_2680/$entry
      -- 
    cp_elements(436) <= cp_elements(25);
    -- CP-element group 437 transition  output  bypass 
    -- predecessors 436 
    -- successors 440 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_2654_to_assign_stmt_2680/AND_u32_u32_2653_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_2654_to_assign_stmt_2680/AND_u32_u32_2653_Update/$entry
      -- 	branch_block_stmt_2042/assign_stmt_2654_to_assign_stmt_2680/AND_u32_u32_2653_Update/cr
      -- 
    cp_elements(437) <= cp_elements(436);
    cr_12089_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(437), ack => AND_u32_u32_2653_inst_req_1); -- 
    -- CP-element group 438 transition  output  bypass 
    -- predecessors 436 
    -- successors 439 
    -- members (7) 
      -- 	branch_block_stmt_2042/assign_stmt_2654_to_assign_stmt_2680/AND_u32_u32_2653_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_2654_to_assign_stmt_2680/R_tempx_x0x_xlcssax_xix_xi50_2650_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_2654_to_assign_stmt_2680/R_tempx_x0x_xlcssax_xix_xi50_2650_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2654_to_assign_stmt_2680/R_tempx_x0x_xlcssax_xix_xi50_2650_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_2654_to_assign_stmt_2680/R_tempx_x0x_xlcssax_xix_xi50_2650_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2654_to_assign_stmt_2680/AND_u32_u32_2653_Sample/$entry
      -- 	branch_block_stmt_2042/assign_stmt_2654_to_assign_stmt_2680/AND_u32_u32_2653_Sample/rr
      -- 
    cp_elements(438) <= cp_elements(436);
    rr_12084_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(438), ack => AND_u32_u32_2653_inst_req_0); -- 
    -- CP-element group 439 transition  input  bypass 
    -- predecessors 438 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_2654_to_assign_stmt_2680/AND_u32_u32_2653_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2654_to_assign_stmt_2680/AND_u32_u32_2653_Sample/$exit
      -- 	branch_block_stmt_2042/assign_stmt_2654_to_assign_stmt_2680/AND_u32_u32_2653_Sample/ra
      -- 
    ra_12085_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => AND_u32_u32_2653_inst_ack_0, ack => cp_elements(439)); -- 
    -- CP-element group 440 transition  input  bypass 
    -- predecessors 437 
    -- successors 448 
    -- members (7) 
      -- 	branch_block_stmt_2042/assign_stmt_2654_to_assign_stmt_2680/AND_u32_u32_2653_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2654_to_assign_stmt_2680/AND_u32_u32_2653_Update/$exit
      -- 	branch_block_stmt_2042/assign_stmt_2654_to_assign_stmt_2680/AND_u32_u32_2653_Update/ca
      -- 	branch_block_stmt_2042/assign_stmt_2654_to_assign_stmt_2680/R_iNsTr_177_2668_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_2654_to_assign_stmt_2680/R_iNsTr_177_2668_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2654_to_assign_stmt_2680/R_iNsTr_177_2668_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_2654_to_assign_stmt_2680/R_iNsTr_177_2668_update_completed_
      -- 
    ca_12090_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => AND_u32_u32_2653_inst_ack_1, ack => cp_elements(440)); -- 
    -- CP-element group 441 transition  output  bypass 
    -- predecessors 436 
    -- successors 444 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_2654_to_assign_stmt_2680/SHL_u32_u32_2659_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_2654_to_assign_stmt_2680/SHL_u32_u32_2659_Update/$entry
      -- 	branch_block_stmt_2042/assign_stmt_2654_to_assign_stmt_2680/SHL_u32_u32_2659_Update/cr
      -- 
    cp_elements(441) <= cp_elements(436);
    cr_12107_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(441), ack => SHL_u32_u32_2659_inst_req_1); -- 
    -- CP-element group 442 transition  output  bypass 
    -- predecessors 436 
    -- successors 443 
    -- members (7) 
      -- 	branch_block_stmt_2042/assign_stmt_2654_to_assign_stmt_2680/SHL_u32_u32_2659_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_2654_to_assign_stmt_2680/R_expx_x0x_xlcssax_xix_xi49_2656_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_2654_to_assign_stmt_2680/R_expx_x0x_xlcssax_xix_xi49_2656_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2654_to_assign_stmt_2680/R_expx_x0x_xlcssax_xix_xi49_2656_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_2654_to_assign_stmt_2680/R_expx_x0x_xlcssax_xix_xi49_2656_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2654_to_assign_stmt_2680/SHL_u32_u32_2659_Sample/$entry
      -- 	branch_block_stmt_2042/assign_stmt_2654_to_assign_stmt_2680/SHL_u32_u32_2659_Sample/rr
      -- 
    cp_elements(442) <= cp_elements(436);
    rr_12102_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(442), ack => SHL_u32_u32_2659_inst_req_0); -- 
    -- CP-element group 443 transition  input  bypass 
    -- predecessors 442 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_2654_to_assign_stmt_2680/SHL_u32_u32_2659_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2654_to_assign_stmt_2680/SHL_u32_u32_2659_Sample/$exit
      -- 	branch_block_stmt_2042/assign_stmt_2654_to_assign_stmt_2680/SHL_u32_u32_2659_Sample/ra
      -- 
    ra_12103_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => SHL_u32_u32_2659_inst_ack_0, ack => cp_elements(443)); -- 
    -- CP-element group 444 transition  input  output  bypass 
    -- predecessors 441 
    -- successors 446 
    -- members (10) 
      -- 	branch_block_stmt_2042/assign_stmt_2654_to_assign_stmt_2680/SHL_u32_u32_2659_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2654_to_assign_stmt_2680/SHL_u32_u32_2659_Update/$exit
      -- 	branch_block_stmt_2042/assign_stmt_2654_to_assign_stmt_2680/SHL_u32_u32_2659_Update/ca
      -- 	branch_block_stmt_2042/assign_stmt_2654_to_assign_stmt_2680/ADD_u32_u32_2665_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_2654_to_assign_stmt_2680/R_iNsTr_178_2662_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_2654_to_assign_stmt_2680/R_iNsTr_178_2662_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2654_to_assign_stmt_2680/R_iNsTr_178_2662_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_2654_to_assign_stmt_2680/R_iNsTr_178_2662_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2654_to_assign_stmt_2680/ADD_u32_u32_2665_Sample/$entry
      -- 	branch_block_stmt_2042/assign_stmt_2654_to_assign_stmt_2680/ADD_u32_u32_2665_Sample/rr
      -- 
    ca_12108_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => SHL_u32_u32_2659_inst_ack_1, ack => cp_elements(444)); -- 
    rr_12120_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(444), ack => ADD_u32_u32_2665_inst_req_0); -- 
    -- CP-element group 445 transition  output  bypass 
    -- predecessors 436 
    -- successors 447 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_2654_to_assign_stmt_2680/ADD_u32_u32_2665_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_2654_to_assign_stmt_2680/ADD_u32_u32_2665_Update/$entry
      -- 	branch_block_stmt_2042/assign_stmt_2654_to_assign_stmt_2680/ADD_u32_u32_2665_Update/cr
      -- 
    cp_elements(445) <= cp_elements(436);
    cr_12125_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(445), ack => ADD_u32_u32_2665_inst_req_1); -- 
    -- CP-element group 446 transition  input  bypass 
    -- predecessors 444 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_2654_to_assign_stmt_2680/ADD_u32_u32_2665_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2654_to_assign_stmt_2680/ADD_u32_u32_2665_Sample/$exit
      -- 	branch_block_stmt_2042/assign_stmt_2654_to_assign_stmt_2680/ADD_u32_u32_2665_Sample/ra
      -- 
    ra_12121_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u32_u32_2665_inst_ack_0, ack => cp_elements(446)); -- 
    -- CP-element group 447 transition  input  bypass 
    -- predecessors 445 
    -- successors 453 
    -- members (7) 
      -- 	branch_block_stmt_2042/assign_stmt_2654_to_assign_stmt_2680/ADD_u32_u32_2665_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2654_to_assign_stmt_2680/ADD_u32_u32_2665_Update/$exit
      -- 	branch_block_stmt_2042/assign_stmt_2654_to_assign_stmt_2680/ADD_u32_u32_2665_Update/ca
      -- 	branch_block_stmt_2042/assign_stmt_2654_to_assign_stmt_2680/R_iNsTr_179_2674_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_2654_to_assign_stmt_2680/R_iNsTr_179_2674_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2654_to_assign_stmt_2680/R_iNsTr_179_2674_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_2654_to_assign_stmt_2680/R_iNsTr_179_2674_update_completed_
      -- 
    ca_12126_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u32_u32_2665_inst_ack_1, ack => cp_elements(447)); -- 
    -- CP-element group 448 join  transition  output  bypass 
    -- predecessors 440 450 
    -- successors 451 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_2654_to_assign_stmt_2680/OR_u32_u32_2670_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_2654_to_assign_stmt_2680/OR_u32_u32_2670_Sample/$entry
      -- 	branch_block_stmt_2042/assign_stmt_2654_to_assign_stmt_2680/OR_u32_u32_2670_Sample/rr
      -- 
    cp_element_group_448: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 20) := "cp_element_group_448"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(440) & cp_elements(450);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(448), clk => clk, reset => reset); --
    end block;
    rr_12142_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(448), ack => OR_u32_u32_2670_inst_req_0); -- 
    -- CP-element group 449 transition  output  bypass 
    -- predecessors 436 
    -- successors 452 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_2654_to_assign_stmt_2680/OR_u32_u32_2670_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_2654_to_assign_stmt_2680/OR_u32_u32_2670_Update/$entry
      -- 	branch_block_stmt_2042/assign_stmt_2654_to_assign_stmt_2680/OR_u32_u32_2670_Update/cr
      -- 
    cp_elements(449) <= cp_elements(436);
    cr_12147_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(449), ack => OR_u32_u32_2670_inst_req_1); -- 
    -- CP-element group 450 transition  bypass 
    -- predecessors 436 
    -- successors 448 
    -- members (4) 
      -- 	branch_block_stmt_2042/assign_stmt_2654_to_assign_stmt_2680/R_iNsTr_140_2669_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_2654_to_assign_stmt_2680/R_iNsTr_140_2669_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2654_to_assign_stmt_2680/R_iNsTr_140_2669_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_2654_to_assign_stmt_2680/R_iNsTr_140_2669_update_completed_
      -- 
    cp_elements(450) <= cp_elements(436);
    -- CP-element group 451 transition  input  bypass 
    -- predecessors 448 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_2654_to_assign_stmt_2680/OR_u32_u32_2670_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2654_to_assign_stmt_2680/OR_u32_u32_2670_Sample/$exit
      -- 	branch_block_stmt_2042/assign_stmt_2654_to_assign_stmt_2680/OR_u32_u32_2670_Sample/ra
      -- 
    ra_12143_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => OR_u32_u32_2670_inst_ack_0, ack => cp_elements(451)); -- 
    -- CP-element group 452 transition  input  bypass 
    -- predecessors 449 
    -- successors 453 
    -- members (7) 
      -- 	branch_block_stmt_2042/assign_stmt_2654_to_assign_stmt_2680/OR_u32_u32_2670_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2654_to_assign_stmt_2680/OR_u32_u32_2670_Update/$exit
      -- 	branch_block_stmt_2042/assign_stmt_2654_to_assign_stmt_2680/OR_u32_u32_2670_Update/ca
      -- 	branch_block_stmt_2042/assign_stmt_2654_to_assign_stmt_2680/R_iNsTr_180_2673_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_2654_to_assign_stmt_2680/R_iNsTr_180_2673_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2654_to_assign_stmt_2680/R_iNsTr_180_2673_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_2654_to_assign_stmt_2680/R_iNsTr_180_2673_update_completed_
      -- 
    ca_12148_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => OR_u32_u32_2670_inst_ack_1, ack => cp_elements(452)); -- 
    -- CP-element group 453 join  transition  output  bypass 
    -- predecessors 447 452 
    -- successors 455 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_2654_to_assign_stmt_2680/OR_u32_u32_2675_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_2654_to_assign_stmt_2680/OR_u32_u32_2675_Sample/$entry
      -- 	branch_block_stmt_2042/assign_stmt_2654_to_assign_stmt_2680/OR_u32_u32_2675_Sample/rr
      -- 
    cp_element_group_453: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 20) := "cp_element_group_453"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(447) & cp_elements(452);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(453), clk => clk, reset => reset); --
    end block;
    rr_12164_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(453), ack => OR_u32_u32_2675_inst_req_0); -- 
    -- CP-element group 454 transition  output  bypass 
    -- predecessors 436 
    -- successors 456 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_2654_to_assign_stmt_2680/OR_u32_u32_2675_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_2654_to_assign_stmt_2680/OR_u32_u32_2675_Update/$entry
      -- 	branch_block_stmt_2042/assign_stmt_2654_to_assign_stmt_2680/OR_u32_u32_2675_Update/cr
      -- 
    cp_elements(454) <= cp_elements(436);
    cr_12169_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(454), ack => OR_u32_u32_2675_inst_req_1); -- 
    -- CP-element group 455 transition  input  bypass 
    -- predecessors 453 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_2654_to_assign_stmt_2680/OR_u32_u32_2675_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2654_to_assign_stmt_2680/OR_u32_u32_2675_Sample/$exit
      -- 	branch_block_stmt_2042/assign_stmt_2654_to_assign_stmt_2680/OR_u32_u32_2675_Sample/ra
      -- 
    ra_12165_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => OR_u32_u32_2675_inst_ack_0, ack => cp_elements(455)); -- 
    -- CP-element group 456 transition  input  output  bypass 
    -- predecessors 454 
    -- successors 458 
    -- members (10) 
      -- 	branch_block_stmt_2042/assign_stmt_2654_to_assign_stmt_2680/type_cast_2679_Sample/rr
      -- 	branch_block_stmt_2042/assign_stmt_2654_to_assign_stmt_2680/type_cast_2679_Sample/$entry
      -- 	branch_block_stmt_2042/assign_stmt_2654_to_assign_stmt_2680/R_iNsTr_181_2678_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2654_to_assign_stmt_2680/OR_u32_u32_2675_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2654_to_assign_stmt_2680/OR_u32_u32_2675_Update/$exit
      -- 	branch_block_stmt_2042/assign_stmt_2654_to_assign_stmt_2680/OR_u32_u32_2675_Update/ca
      -- 	branch_block_stmt_2042/assign_stmt_2654_to_assign_stmt_2680/type_cast_2679_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_2654_to_assign_stmt_2680/R_iNsTr_181_2678_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_2654_to_assign_stmt_2680/R_iNsTr_181_2678_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2654_to_assign_stmt_2680/R_iNsTr_181_2678_update_start_
      -- 
    ca_12170_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => OR_u32_u32_2675_inst_ack_1, ack => cp_elements(456)); -- 
    rr_12182_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(456), ack => type_cast_2679_inst_req_0); -- 
    -- CP-element group 457 transition  output  bypass 
    -- predecessors 436 
    -- successors 459 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_2654_to_assign_stmt_2680/type_cast_2679_Update/cr
      -- 	branch_block_stmt_2042/assign_stmt_2654_to_assign_stmt_2680/type_cast_2679_Update/$entry
      -- 	branch_block_stmt_2042/assign_stmt_2654_to_assign_stmt_2680/type_cast_2679_update_start_
      -- 
    cp_elements(457) <= cp_elements(436);
    cr_12187_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(457), ack => type_cast_2679_inst_req_1); -- 
    -- CP-element group 458 transition  input  bypass 
    -- predecessors 456 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_2654_to_assign_stmt_2680/type_cast_2679_Sample/ra
      -- 	branch_block_stmt_2042/assign_stmt_2654_to_assign_stmt_2680/type_cast_2679_Sample/$exit
      -- 	branch_block_stmt_2042/assign_stmt_2654_to_assign_stmt_2680/type_cast_2679_sample_completed_
      -- 
    ra_12183_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2679_inst_ack_0, ack => cp_elements(458)); -- 
    -- CP-element group 459 fork  transition  place  input  bypass 
    -- predecessors 457 
    -- successors 1654 1656 
    -- members (11) 
      -- 	branch_block_stmt_2042/assign_stmt_2654_to_assign_stmt_2680__exit__
      -- 	branch_block_stmt_2042/xx_xcritedgex_xix_xi52_rotor_flux_calcx_xexit
      -- 	branch_block_stmt_2042/assign_stmt_2654_to_assign_stmt_2680/type_cast_2679_Update/ca
      -- 	branch_block_stmt_2042/assign_stmt_2654_to_assign_stmt_2680/type_cast_2679_Update/$exit
      -- 	branch_block_stmt_2042/assign_stmt_2654_to_assign_stmt_2680/$exit
      -- 	branch_block_stmt_2042/assign_stmt_2654_to_assign_stmt_2680/type_cast_2679_update_completed_
      -- 	branch_block_stmt_2042/xx_xcritedgex_xix_xi52_rotor_flux_calcx_xexit_PhiReq/phi_stmt_2683/phi_stmt_2683_sources/type_cast_2686/SplitProtocol/$entry
      -- 	branch_block_stmt_2042/xx_xcritedgex_xix_xi52_rotor_flux_calcx_xexit_PhiReq/$entry
      -- 	branch_block_stmt_2042/xx_xcritedgex_xix_xi52_rotor_flux_calcx_xexit_PhiReq/phi_stmt_2683/$entry
      -- 	branch_block_stmt_2042/xx_xcritedgex_xix_xi52_rotor_flux_calcx_xexit_PhiReq/phi_stmt_2683/phi_stmt_2683_sources/$entry
      -- 	branch_block_stmt_2042/xx_xcritedgex_xix_xi52_rotor_flux_calcx_xexit_PhiReq/phi_stmt_2683/phi_stmt_2683_sources/type_cast_2686/$entry
      -- 
    ca_12188_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2679_inst_ack_1, ack => cp_elements(459)); -- 
    -- CP-element group 460 fork  transition  bypass 
    -- predecessors 1661 
    -- successors 461 462 465 466 469 473 476 
    -- members (1) 
      -- 	branch_block_stmt_2042/assign_stmt_2696_to_assign_stmt_2716/$entry
      -- 
    cp_elements(460) <= cp_elements(1661);
    -- CP-element group 461 transition  output  bypass 
    -- predecessors 460 
    -- successors 464 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_2696_to_assign_stmt_2716/MUL_f32_f32_2695_Update/$entry
      -- 	branch_block_stmt_2042/assign_stmt_2696_to_assign_stmt_2716/MUL_f32_f32_2695_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_2696_to_assign_stmt_2716/MUL_f32_f32_2695_Update/cr
      -- 
    cp_elements(461) <= cp_elements(460);
    cr_12208_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(461), ack => MUL_f32_f32_2695_inst_req_1); -- 
    -- CP-element group 462 transition  output  bypass 
    -- predecessors 460 
    -- successors 463 
    -- members (7) 
      -- 	branch_block_stmt_2042/assign_stmt_2696_to_assign_stmt_2716/R_iNsTr_4_2692_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_2696_to_assign_stmt_2716/R_iNsTr_4_2692_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2696_to_assign_stmt_2716/MUL_f32_f32_2695_Sample/$entry
      -- 	branch_block_stmt_2042/assign_stmt_2696_to_assign_stmt_2716/MUL_f32_f32_2695_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_2696_to_assign_stmt_2716/MUL_f32_f32_2695_Sample/rr
      -- 	branch_block_stmt_2042/assign_stmt_2696_to_assign_stmt_2716/R_iNsTr_4_2692_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2696_to_assign_stmt_2716/R_iNsTr_4_2692_sample_start_
      -- 
    cp_elements(462) <= cp_elements(460);
    rr_12203_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(462), ack => MUL_f32_f32_2695_inst_req_0); -- 
    -- CP-element group 463 transition  input  bypass 
    -- predecessors 462 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_2696_to_assign_stmt_2716/MUL_f32_f32_2695_Sample/ra
      -- 	branch_block_stmt_2042/assign_stmt_2696_to_assign_stmt_2716/MUL_f32_f32_2695_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2696_to_assign_stmt_2716/MUL_f32_f32_2695_Sample/$exit
      -- 
    ra_12204_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => MUL_f32_f32_2695_inst_ack_0, ack => cp_elements(463)); -- 
    -- CP-element group 464 fork  transition  input  bypass 
    -- predecessors 461 
    -- successors 470 477 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_2696_to_assign_stmt_2716/MUL_f32_f32_2695_Update/ca
      -- 	branch_block_stmt_2042/assign_stmt_2696_to_assign_stmt_2716/MUL_f32_f32_2695_Update/$exit
      -- 	branch_block_stmt_2042/assign_stmt_2696_to_assign_stmt_2716/MUL_f32_f32_2695_update_completed_
      -- 
    ca_12209_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => MUL_f32_f32_2695_inst_ack_1, ack => cp_elements(464)); -- 
    -- CP-element group 465 transition  output  bypass 
    -- predecessors 460 
    -- successors 468 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_2696_to_assign_stmt_2716/MUL_f32_f32_2701_Update/cr
      -- 	branch_block_stmt_2042/assign_stmt_2696_to_assign_stmt_2716/MUL_f32_f32_2701_Update/$entry
      -- 	branch_block_stmt_2042/assign_stmt_2696_to_assign_stmt_2716/MUL_f32_f32_2701_update_start_
      -- 
    cp_elements(465) <= cp_elements(460);
    cr_12226_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(465), ack => MUL_f32_f32_2701_inst_req_1); -- 
    -- CP-element group 466 transition  output  bypass 
    -- predecessors 460 
    -- successors 467 
    -- members (7) 
      -- 	branch_block_stmt_2042/assign_stmt_2696_to_assign_stmt_2716/MUL_f32_f32_2701_Sample/rr
      -- 	branch_block_stmt_2042/assign_stmt_2696_to_assign_stmt_2716/MUL_f32_f32_2701_Sample/$entry
      -- 	branch_block_stmt_2042/assign_stmt_2696_to_assign_stmt_2716/R_iNsTr_42_2698_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2696_to_assign_stmt_2716/R_iNsTr_42_2698_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_2696_to_assign_stmt_2716/R_iNsTr_42_2698_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2696_to_assign_stmt_2716/R_iNsTr_42_2698_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_2696_to_assign_stmt_2716/MUL_f32_f32_2701_sample_start_
      -- 
    cp_elements(466) <= cp_elements(460);
    rr_12221_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(466), ack => MUL_f32_f32_2701_inst_req_0); -- 
    -- CP-element group 467 transition  input  bypass 
    -- predecessors 466 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_2696_to_assign_stmt_2716/MUL_f32_f32_2701_Sample/ra
      -- 	branch_block_stmt_2042/assign_stmt_2696_to_assign_stmt_2716/MUL_f32_f32_2701_Sample/$exit
      -- 	branch_block_stmt_2042/assign_stmt_2696_to_assign_stmt_2716/MUL_f32_f32_2701_sample_completed_
      -- 
    ra_12222_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => MUL_f32_f32_2701_inst_ack_0, ack => cp_elements(467)); -- 
    -- CP-element group 468 transition  input  output  bypass 
    -- predecessors 465 
    -- successors 474 
    -- members (10) 
      -- 	branch_block_stmt_2042/assign_stmt_2696_to_assign_stmt_2716/type_cast_2709_Sample/rr
      -- 	branch_block_stmt_2042/assign_stmt_2696_to_assign_stmt_2716/type_cast_2709_Sample/$entry
      -- 	branch_block_stmt_2042/assign_stmt_2696_to_assign_stmt_2716/R_iNsTr_44_2708_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2696_to_assign_stmt_2716/R_iNsTr_44_2708_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_2696_to_assign_stmt_2716/R_iNsTr_44_2708_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2696_to_assign_stmt_2716/R_iNsTr_44_2708_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_2696_to_assign_stmt_2716/type_cast_2709_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_2696_to_assign_stmt_2716/MUL_f32_f32_2701_Update/ca
      -- 	branch_block_stmt_2042/assign_stmt_2696_to_assign_stmt_2716/MUL_f32_f32_2701_Update/$exit
      -- 	branch_block_stmt_2042/assign_stmt_2696_to_assign_stmt_2716/MUL_f32_f32_2701_update_completed_
      -- 
    ca_12227_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => MUL_f32_f32_2701_inst_ack_1, ack => cp_elements(468)); -- 
    rr_12257_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(468), ack => type_cast_2709_inst_req_0); -- 
    -- CP-element group 469 transition  output  bypass 
    -- predecessors 460 
    -- successors 472 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_2696_to_assign_stmt_2716/type_cast_2705_Update/cr
      -- 	branch_block_stmt_2042/assign_stmt_2696_to_assign_stmt_2716/type_cast_2705_Update/$entry
      -- 	branch_block_stmt_2042/assign_stmt_2696_to_assign_stmt_2716/type_cast_2705_update_start_
      -- 
    cp_elements(469) <= cp_elements(460);
    cr_12244_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(469), ack => type_cast_2705_inst_req_1); -- 
    -- CP-element group 470 transition  output  bypass 
    -- predecessors 464 
    -- successors 471 
    -- members (7) 
      -- 	branch_block_stmt_2042/assign_stmt_2696_to_assign_stmt_2716/type_cast_2705_Sample/rr
      -- 	branch_block_stmt_2042/assign_stmt_2696_to_assign_stmt_2716/type_cast_2705_Sample/$entry
      -- 	branch_block_stmt_2042/assign_stmt_2696_to_assign_stmt_2716/R_iNsTr_43_2704_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2696_to_assign_stmt_2716/R_iNsTr_43_2704_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_2696_to_assign_stmt_2716/R_iNsTr_43_2704_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2696_to_assign_stmt_2716/R_iNsTr_43_2704_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_2696_to_assign_stmt_2716/type_cast_2705_sample_start_
      -- 
    cp_elements(470) <= cp_elements(464);
    rr_12239_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(470), ack => type_cast_2705_inst_req_0); -- 
    -- CP-element group 471 transition  input  bypass 
    -- predecessors 470 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_2696_to_assign_stmt_2716/type_cast_2705_Sample/ra
      -- 	branch_block_stmt_2042/assign_stmt_2696_to_assign_stmt_2716/type_cast_2705_Sample/$exit
      -- 	branch_block_stmt_2042/assign_stmt_2696_to_assign_stmt_2716/type_cast_2705_sample_completed_
      -- 
    ra_12240_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2705_inst_ack_0, ack => cp_elements(471)); -- 
    -- CP-element group 472 transition  input  bypass 
    -- predecessors 469 
    -- successors 480 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_2696_to_assign_stmt_2716/type_cast_2705_Update/ca
      -- 	branch_block_stmt_2042/assign_stmt_2696_to_assign_stmt_2716/type_cast_2705_Update/$exit
      -- 	branch_block_stmt_2042/assign_stmt_2696_to_assign_stmt_2716/type_cast_2705_update_completed_
      -- 
    ca_12245_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2705_inst_ack_1, ack => cp_elements(472)); -- 
    -- CP-element group 473 transition  output  bypass 
    -- predecessors 460 
    -- successors 475 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_2696_to_assign_stmt_2716/type_cast_2709_Update/cr
      -- 	branch_block_stmt_2042/assign_stmt_2696_to_assign_stmt_2716/type_cast_2709_Update/$entry
      -- 	branch_block_stmt_2042/assign_stmt_2696_to_assign_stmt_2716/type_cast_2709_update_start_
      -- 
    cp_elements(473) <= cp_elements(460);
    cr_12262_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(473), ack => type_cast_2709_inst_req_1); -- 
    -- CP-element group 474 transition  input  bypass 
    -- predecessors 468 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_2696_to_assign_stmt_2716/type_cast_2709_Sample/ra
      -- 	branch_block_stmt_2042/assign_stmt_2696_to_assign_stmt_2716/type_cast_2709_Sample/$exit
      -- 	branch_block_stmt_2042/assign_stmt_2696_to_assign_stmt_2716/type_cast_2709_sample_completed_
      -- 
    ra_12258_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2709_inst_ack_0, ack => cp_elements(474)); -- 
    -- CP-element group 475 transition  input  bypass 
    -- predecessors 473 
    -- successors 480 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_2696_to_assign_stmt_2716/type_cast_2709_Update/ca
      -- 	branch_block_stmt_2042/assign_stmt_2696_to_assign_stmt_2716/type_cast_2709_Update/$exit
      -- 	branch_block_stmt_2042/assign_stmt_2696_to_assign_stmt_2716/type_cast_2709_update_completed_
      -- 
    ca_12263_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2709_inst_ack_1, ack => cp_elements(475)); -- 
    -- CP-element group 476 transition  output  bypass 
    -- predecessors 460 
    -- successors 479 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_2696_to_assign_stmt_2716/EQ_f32_u1_2715_Update/$entry
      -- 	branch_block_stmt_2042/assign_stmt_2696_to_assign_stmt_2716/EQ_f32_u1_2715_Update/cr
      -- 	branch_block_stmt_2042/assign_stmt_2696_to_assign_stmt_2716/EQ_f32_u1_2715_update_start_
      -- 
    cp_elements(476) <= cp_elements(460);
    cr_12280_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(476), ack => EQ_f32_u1_2715_inst_req_1); -- 
    -- CP-element group 477 transition  output  bypass 
    -- predecessors 464 
    -- successors 478 
    -- members (7) 
      -- 	branch_block_stmt_2042/assign_stmt_2696_to_assign_stmt_2716/R_iNsTr_43_2712_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2696_to_assign_stmt_2716/R_iNsTr_43_2712_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_2696_to_assign_stmt_2716/R_iNsTr_43_2712_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2696_to_assign_stmt_2716/EQ_f32_u1_2715_Sample/$entry
      -- 	branch_block_stmt_2042/assign_stmt_2696_to_assign_stmt_2716/EQ_f32_u1_2715_Sample/rr
      -- 	branch_block_stmt_2042/assign_stmt_2696_to_assign_stmt_2716/R_iNsTr_43_2712_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_2696_to_assign_stmt_2716/EQ_f32_u1_2715_sample_start_
      -- 
    cp_elements(477) <= cp_elements(464);
    rr_12275_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(477), ack => EQ_f32_u1_2715_inst_req_0); -- 
    -- CP-element group 478 transition  input  bypass 
    -- predecessors 477 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_2696_to_assign_stmt_2716/EQ_f32_u1_2715_Sample/$exit
      -- 	branch_block_stmt_2042/assign_stmt_2696_to_assign_stmt_2716/EQ_f32_u1_2715_Sample/ra
      -- 	branch_block_stmt_2042/assign_stmt_2696_to_assign_stmt_2716/EQ_f32_u1_2715_sample_completed_
      -- 
    ra_12276_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_f32_u1_2715_inst_ack_0, ack => cp_elements(478)); -- 
    -- CP-element group 479 transition  input  bypass 
    -- predecessors 476 
    -- successors 480 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_2696_to_assign_stmt_2716/EQ_f32_u1_2715_Update/$exit
      -- 	branch_block_stmt_2042/assign_stmt_2696_to_assign_stmt_2716/EQ_f32_u1_2715_Update/ca
      -- 	branch_block_stmt_2042/assign_stmt_2696_to_assign_stmt_2716/EQ_f32_u1_2715_update_completed_
      -- 
    ca_12281_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_f32_u1_2715_inst_ack_1, ack => cp_elements(479)); -- 
    -- CP-element group 480 join  transition  bypass 
    -- predecessors 472 475 479 
    -- successors 26 
    -- members (1) 
      -- 	branch_block_stmt_2042/assign_stmt_2696_to_assign_stmt_2716/$exit
      -- 
    cp_element_group_480: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 20) := "cp_element_group_480"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= cp_elements(472) & cp_elements(475) & cp_elements(479);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(480), clk => clk, reset => reset); --
    end block;
    -- CP-element group 481 transition  place  dead  bypass 
    -- predecessors 26 
    -- successors 27 
    -- members (8) 
      -- 	branch_block_stmt_2042/merge_stmt_2723__entry__
      -- 	branch_block_stmt_2042/if_stmt_2717__exit__
      -- 	branch_block_stmt_2042/if_stmt_2717_dead_link/$exit
      -- 	branch_block_stmt_2042/if_stmt_2717_dead_link/$entry
      -- 	branch_block_stmt_2042/if_stmt_2717_dead_link/dead_transition
      -- 	branch_block_stmt_2042/merge_stmt_2723_dead_link/dead_transition
      -- 	branch_block_stmt_2042/merge_stmt_2723_dead_link/$exit
      -- 	branch_block_stmt_2042/merge_stmt_2723_dead_link/$entry
      -- 
    cp_elements(481) <= false;
    -- CP-element group 482 transition  output  bypass 
    -- predecessors 26 
    -- successors 483 
    -- members (3) 
      -- 	branch_block_stmt_2042/if_stmt_2717_eval_test/$entry
      -- 	branch_block_stmt_2042/if_stmt_2717_eval_test/branch_req
      -- 	branch_block_stmt_2042/if_stmt_2717_eval_test/$exit
      -- 
    cp_elements(482) <= cp_elements(26);
    branch_req_12289_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(482), ack => if_stmt_2717_branch_req_0); -- 
    -- CP-element group 483 branch  place  bypass 
    -- predecessors 482 
    -- successors 484 486 
    -- members (1) 
      -- 	branch_block_stmt_2042/R_iNsTr_45_2718_place
      -- 
    cp_elements(483) <= cp_elements(482);
    -- CP-element group 484 transition  bypass 
    -- predecessors 483 
    -- successors 485 
    -- members (1) 
      -- 	branch_block_stmt_2042/if_stmt_2717_if_link/$entry
      -- 
    cp_elements(484) <= cp_elements(483);
    -- CP-element group 485 fork  transition  place  input  bypass 
    -- predecessors 484 
    -- successors 1971 1972 
    -- members (8) 
      -- 	branch_block_stmt_2042/if_stmt_2717_if_link/if_choice_transition
      -- 	branch_block_stmt_2042/if_stmt_2717_if_link/$exit
      -- 	branch_block_stmt_2042/rotor_flux_calcx_xexit_omega_calcx_xexit
      -- 	branch_block_stmt_2042/rotor_flux_calcx_xexit_omega_calcx_xexit_PhiReq/$entry
      -- 	branch_block_stmt_2042/rotor_flux_calcx_xexit_omega_calcx_xexit_PhiReq/phi_stmt_3122/$entry
      -- 	branch_block_stmt_2042/rotor_flux_calcx_xexit_omega_calcx_xexit_PhiReq/phi_stmt_3122/phi_stmt_3122_sources/$entry
      -- 	branch_block_stmt_2042/rotor_flux_calcx_xexit_omega_calcx_xexit_PhiReq/phi_stmt_3122/phi_stmt_3122_sources/type_cast_3125/$entry
      -- 	branch_block_stmt_2042/rotor_flux_calcx_xexit_omega_calcx_xexit_PhiReq/phi_stmt_3122/phi_stmt_3122_sources/type_cast_3125/SplitProtocol/$entry
      -- 
    if_choice_transition_12294_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2717_branch_ack_1, ack => cp_elements(485)); -- 
    -- CP-element group 486 transition  bypass 
    -- predecessors 483 
    -- successors 487 
    -- members (1) 
      -- 	branch_block_stmt_2042/if_stmt_2717_else_link/$entry
      -- 
    cp_elements(486) <= cp_elements(483);
    -- CP-element group 487 transition  place  input  bypass 
    -- predecessors 486 
    -- successors 27 
    -- members (9) 
      -- 	branch_block_stmt_2042/if_stmt_2717_else_link/else_choice_transition
      -- 	branch_block_stmt_2042/if_stmt_2717_else_link/$exit
      -- 	branch_block_stmt_2042/rotor_flux_calcx_xexit_bb_26
      -- 	branch_block_stmt_2042/merge_stmt_2723_PhiAck/$entry
      -- 	branch_block_stmt_2042/merge_stmt_2723_PhiAck/$exit
      -- 	branch_block_stmt_2042/rotor_flux_calcx_xexit_bb_26_PhiReq/$exit
      -- 	branch_block_stmt_2042/rotor_flux_calcx_xexit_bb_26_PhiReq/$entry
      -- 	branch_block_stmt_2042/merge_stmt_2723_PhiAck/dummy
      -- 	branch_block_stmt_2042/merge_stmt_2723_PhiReqMerge
      -- 
    else_choice_transition_12298_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2717_branch_ack_0, ack => cp_elements(487)); -- 
    -- CP-element group 488 fork  transition  bypass 
    -- predecessors 27 
    -- successors 489 490 493 496 497 500 503 504 507 510 513 514 517 520 524 525 526 529 533 
    -- members (1) 
      -- 	branch_block_stmt_2042/assign_stmt_2729_to_assign_stmt_2799/$entry
      -- 
    cp_elements(488) <= cp_elements(27);
    -- CP-element group 489 transition  output  bypass 
    -- predecessors 488 
    -- successors 492 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_2729_to_assign_stmt_2799/LSHR_u32_u32_2728_Update/$entry
      -- 	branch_block_stmt_2042/assign_stmt_2729_to_assign_stmt_2799/LSHR_u32_u32_2728_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_2729_to_assign_stmt_2799/LSHR_u32_u32_2728_Update/cr
      -- 
    cp_elements(489) <= cp_elements(488);
    cr_12320_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(489), ack => LSHR_u32_u32_2728_inst_req_1); -- 
    -- CP-element group 490 transition  output  bypass 
    -- predecessors 488 
    -- successors 491 
    -- members (7) 
      -- 	branch_block_stmt_2042/assign_stmt_2729_to_assign_stmt_2799/LSHR_u32_u32_2728_Sample/rr
      -- 	branch_block_stmt_2042/assign_stmt_2729_to_assign_stmt_2799/R_tmp10x_xix_xi1_2725_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_2729_to_assign_stmt_2799/R_tmp10x_xix_xi1_2725_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2729_to_assign_stmt_2799/LSHR_u32_u32_2728_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_2729_to_assign_stmt_2799/LSHR_u32_u32_2728_Sample/$entry
      -- 	branch_block_stmt_2042/assign_stmt_2729_to_assign_stmt_2799/R_tmp10x_xix_xi1_2725_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2729_to_assign_stmt_2799/R_tmp10x_xix_xi1_2725_update_start_
      -- 
    cp_elements(490) <= cp_elements(488);
    rr_12315_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(490), ack => LSHR_u32_u32_2728_inst_req_0); -- 
    -- CP-element group 491 transition  input  bypass 
    -- predecessors 490 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_2729_to_assign_stmt_2799/LSHR_u32_u32_2728_Sample/ra
      -- 	branch_block_stmt_2042/assign_stmt_2729_to_assign_stmt_2799/LSHR_u32_u32_2728_Sample/$exit
      -- 	branch_block_stmt_2042/assign_stmt_2729_to_assign_stmt_2799/LSHR_u32_u32_2728_sample_completed_
      -- 
    ra_12316_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => LSHR_u32_u32_2728_inst_ack_0, ack => cp_elements(491)); -- 
    -- CP-element group 492 transition  input  output  bypass 
    -- predecessors 489 
    -- successors 494 
    -- members (10) 
      -- 	branch_block_stmt_2042/assign_stmt_2729_to_assign_stmt_2799/LSHR_u32_u32_2728_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2729_to_assign_stmt_2799/R_iNsTr_64_2731_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_2729_to_assign_stmt_2799/AND_u32_u32_2734_Sample/$entry
      -- 	branch_block_stmt_2042/assign_stmt_2729_to_assign_stmt_2799/R_iNsTr_64_2731_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2729_to_assign_stmt_2799/AND_u32_u32_2734_Sample/rr
      -- 	branch_block_stmt_2042/assign_stmt_2729_to_assign_stmt_2799/AND_u32_u32_2734_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_2729_to_assign_stmt_2799/LSHR_u32_u32_2728_Update/ca
      -- 	branch_block_stmt_2042/assign_stmt_2729_to_assign_stmt_2799/R_iNsTr_64_2731_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_2729_to_assign_stmt_2799/LSHR_u32_u32_2728_Update/$exit
      -- 	branch_block_stmt_2042/assign_stmt_2729_to_assign_stmt_2799/R_iNsTr_64_2731_sample_completed_
      -- 
    ca_12321_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => LSHR_u32_u32_2728_inst_ack_1, ack => cp_elements(492)); -- 
    rr_12333_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(492), ack => AND_u32_u32_2734_inst_req_0); -- 
    -- CP-element group 493 transition  output  bypass 
    -- predecessors 488 
    -- successors 495 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_2729_to_assign_stmt_2799/AND_u32_u32_2734_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_2729_to_assign_stmt_2799/AND_u32_u32_2734_Update/cr
      -- 	branch_block_stmt_2042/assign_stmt_2729_to_assign_stmt_2799/AND_u32_u32_2734_Update/$entry
      -- 
    cp_elements(493) <= cp_elements(488);
    cr_12338_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(493), ack => AND_u32_u32_2734_inst_req_1); -- 
    -- CP-element group 494 transition  input  bypass 
    -- predecessors 492 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_2729_to_assign_stmt_2799/AND_u32_u32_2734_Sample/$exit
      -- 	branch_block_stmt_2042/assign_stmt_2729_to_assign_stmt_2799/AND_u32_u32_2734_Sample/ra
      -- 	branch_block_stmt_2042/assign_stmt_2729_to_assign_stmt_2799/AND_u32_u32_2734_sample_completed_
      -- 
    ra_12334_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => AND_u32_u32_2734_inst_ack_0, ack => cp_elements(494)); -- 
    -- CP-element group 495 transition  input  bypass 
    -- predecessors 493 
    -- successors 532 
    -- members (7) 
      -- 	branch_block_stmt_2042/assign_stmt_2729_to_assign_stmt_2799/AND_u32_u32_2734_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2729_to_assign_stmt_2799/AND_u32_u32_2734_Update/ca
      -- 	branch_block_stmt_2042/assign_stmt_2729_to_assign_stmt_2799/AND_u32_u32_2734_Update/$exit
      -- 	branch_block_stmt_2042/assign_stmt_2729_to_assign_stmt_2799/R_iNsTr_65_2796_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2729_to_assign_stmt_2799/R_iNsTr_65_2796_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_2729_to_assign_stmt_2799/R_iNsTr_65_2796_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_2729_to_assign_stmt_2799/R_iNsTr_65_2796_update_completed_
      -- 
    ca_12339_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => AND_u32_u32_2734_inst_ack_1, ack => cp_elements(495)); -- 
    -- CP-element group 496 transition  output  bypass 
    -- predecessors 488 
    -- successors 499 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_2729_to_assign_stmt_2799/LSHR_u32_u32_2740_Update/cr
      -- 	branch_block_stmt_2042/assign_stmt_2729_to_assign_stmt_2799/LSHR_u32_u32_2740_Update/$entry
      -- 	branch_block_stmt_2042/assign_stmt_2729_to_assign_stmt_2799/LSHR_u32_u32_2740_update_start_
      -- 
    cp_elements(496) <= cp_elements(488);
    cr_12356_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(496), ack => LSHR_u32_u32_2740_inst_req_1); -- 
    -- CP-element group 497 transition  output  bypass 
    -- predecessors 488 
    -- successors 498 
    -- members (7) 
      -- 	branch_block_stmt_2042/assign_stmt_2729_to_assign_stmt_2799/LSHR_u32_u32_2740_Sample/rr
      -- 	branch_block_stmt_2042/assign_stmt_2729_to_assign_stmt_2799/R_tmp6x_xix_xi2_2737_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_2729_to_assign_stmt_2799/R_tmp6x_xix_xi2_2737_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2729_to_assign_stmt_2799/LSHR_u32_u32_2740_Sample/$entry
      -- 	branch_block_stmt_2042/assign_stmt_2729_to_assign_stmt_2799/R_tmp6x_xix_xi2_2737_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2729_to_assign_stmt_2799/R_tmp6x_xix_xi2_2737_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_2729_to_assign_stmt_2799/LSHR_u32_u32_2740_sample_start_
      -- 
    cp_elements(497) <= cp_elements(488);
    rr_12351_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(497), ack => LSHR_u32_u32_2740_inst_req_0); -- 
    -- CP-element group 498 transition  input  bypass 
    -- predecessors 497 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_2729_to_assign_stmt_2799/LSHR_u32_u32_2740_Sample/ra
      -- 	branch_block_stmt_2042/assign_stmt_2729_to_assign_stmt_2799/LSHR_u32_u32_2740_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2729_to_assign_stmt_2799/LSHR_u32_u32_2740_Sample/$exit
      -- 
    ra_12352_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => LSHR_u32_u32_2740_inst_ack_0, ack => cp_elements(498)); -- 
    -- CP-element group 499 transition  input  output  bypass 
    -- predecessors 496 
    -- successors 501 
    -- members (10) 
      -- 	branch_block_stmt_2042/assign_stmt_2729_to_assign_stmt_2799/LSHR_u32_u32_2740_Update/ca
      -- 	branch_block_stmt_2042/assign_stmt_2729_to_assign_stmt_2799/LSHR_u32_u32_2740_Update/$exit
      -- 	branch_block_stmt_2042/assign_stmt_2729_to_assign_stmt_2799/R_iNsTr_66_2743_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2729_to_assign_stmt_2799/R_iNsTr_66_2743_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_2729_to_assign_stmt_2799/R_iNsTr_66_2743_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2729_to_assign_stmt_2799/LSHR_u32_u32_2740_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2729_to_assign_stmt_2799/AND_u32_u32_2746_Sample/rr
      -- 	branch_block_stmt_2042/assign_stmt_2729_to_assign_stmt_2799/AND_u32_u32_2746_Sample/$entry
      -- 	branch_block_stmt_2042/assign_stmt_2729_to_assign_stmt_2799/R_iNsTr_66_2743_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_2729_to_assign_stmt_2799/AND_u32_u32_2746_sample_start_
      -- 
    ca_12357_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => LSHR_u32_u32_2740_inst_ack_1, ack => cp_elements(499)); -- 
    rr_12369_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(499), ack => AND_u32_u32_2746_inst_req_0); -- 
    -- CP-element group 500 transition  output  bypass 
    -- predecessors 488 
    -- successors 502 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_2729_to_assign_stmt_2799/AND_u32_u32_2746_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_2729_to_assign_stmt_2799/AND_u32_u32_2746_Update/cr
      -- 	branch_block_stmt_2042/assign_stmt_2729_to_assign_stmt_2799/AND_u32_u32_2746_Update/$entry
      -- 
    cp_elements(500) <= cp_elements(488);
    cr_12374_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(500), ack => AND_u32_u32_2746_inst_req_1); -- 
    -- CP-element group 501 transition  input  bypass 
    -- predecessors 499 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_2729_to_assign_stmt_2799/AND_u32_u32_2746_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2729_to_assign_stmt_2799/AND_u32_u32_2746_Sample/ra
      -- 	branch_block_stmt_2042/assign_stmt_2729_to_assign_stmt_2799/AND_u32_u32_2746_Sample/$exit
      -- 
    ra_12370_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => AND_u32_u32_2746_inst_ack_0, ack => cp_elements(501)); -- 
    -- CP-element group 502 transition  input  bypass 
    -- predecessors 500 
    -- successors 532 
    -- members (7) 
      -- 	branch_block_stmt_2042/assign_stmt_2729_to_assign_stmt_2799/AND_u32_u32_2746_Update/ca
      -- 	branch_block_stmt_2042/assign_stmt_2729_to_assign_stmt_2799/AND_u32_u32_2746_Update/$exit
      -- 	branch_block_stmt_2042/assign_stmt_2729_to_assign_stmt_2799/AND_u32_u32_2746_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2729_to_assign_stmt_2799/R_iNsTr_67_2797_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_2729_to_assign_stmt_2799/R_iNsTr_67_2797_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2729_to_assign_stmt_2799/R_iNsTr_67_2797_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_2729_to_assign_stmt_2799/R_iNsTr_67_2797_update_completed_
      -- 
    ca_12375_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => AND_u32_u32_2746_inst_ack_1, ack => cp_elements(502)); -- 
    -- CP-element group 503 transition  output  bypass 
    -- predecessors 488 
    -- successors 506 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_2729_to_assign_stmt_2799/SHL_u32_u32_2752_Update/cr
      -- 	branch_block_stmt_2042/assign_stmt_2729_to_assign_stmt_2799/SHL_u32_u32_2752_Update/$entry
      -- 	branch_block_stmt_2042/assign_stmt_2729_to_assign_stmt_2799/SHL_u32_u32_2752_update_start_
      -- 
    cp_elements(503) <= cp_elements(488);
    cr_12392_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(503), ack => SHL_u32_u32_2752_inst_req_1); -- 
    -- CP-element group 504 transition  output  bypass 
    -- predecessors 488 
    -- successors 505 
    -- members (7) 
      -- 	branch_block_stmt_2042/assign_stmt_2729_to_assign_stmt_2799/SHL_u32_u32_2752_Sample/rr
      -- 	branch_block_stmt_2042/assign_stmt_2729_to_assign_stmt_2799/SHL_u32_u32_2752_Sample/$entry
      -- 	branch_block_stmt_2042/assign_stmt_2729_to_assign_stmt_2799/R_tmp10x_xix_xi1_2749_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2729_to_assign_stmt_2799/R_tmp10x_xix_xi1_2749_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_2729_to_assign_stmt_2799/R_tmp10x_xix_xi1_2749_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2729_to_assign_stmt_2799/R_tmp10x_xix_xi1_2749_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_2729_to_assign_stmt_2799/SHL_u32_u32_2752_sample_start_
      -- 
    cp_elements(504) <= cp_elements(488);
    rr_12387_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(504), ack => SHL_u32_u32_2752_inst_req_0); -- 
    -- CP-element group 505 transition  input  bypass 
    -- predecessors 504 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_2729_to_assign_stmt_2799/SHL_u32_u32_2752_Sample/ra
      -- 	branch_block_stmt_2042/assign_stmt_2729_to_assign_stmt_2799/SHL_u32_u32_2752_Sample/$exit
      -- 	branch_block_stmt_2042/assign_stmt_2729_to_assign_stmt_2799/SHL_u32_u32_2752_sample_completed_
      -- 
    ra_12388_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => SHL_u32_u32_2752_inst_ack_0, ack => cp_elements(505)); -- 
    -- CP-element group 506 transition  input  output  bypass 
    -- predecessors 503 
    -- successors 508 
    -- members (10) 
      -- 	branch_block_stmt_2042/assign_stmt_2729_to_assign_stmt_2799/R_iNsTr_68_2755_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_2729_to_assign_stmt_2799/AND_u32_u32_2758_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_2729_to_assign_stmt_2799/SHL_u32_u32_2752_Update/ca
      -- 	branch_block_stmt_2042/assign_stmt_2729_to_assign_stmt_2799/SHL_u32_u32_2752_Update/$exit
      -- 	branch_block_stmt_2042/assign_stmt_2729_to_assign_stmt_2799/R_iNsTr_68_2755_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2729_to_assign_stmt_2799/AND_u32_u32_2758_Sample/$entry
      -- 	branch_block_stmt_2042/assign_stmt_2729_to_assign_stmt_2799/SHL_u32_u32_2752_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2729_to_assign_stmt_2799/AND_u32_u32_2758_Sample/rr
      -- 	branch_block_stmt_2042/assign_stmt_2729_to_assign_stmt_2799/R_iNsTr_68_2755_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2729_to_assign_stmt_2799/R_iNsTr_68_2755_update_start_
      -- 
    ca_12393_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => SHL_u32_u32_2752_inst_ack_1, ack => cp_elements(506)); -- 
    rr_12405_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(506), ack => AND_u32_u32_2758_inst_req_0); -- 
    -- CP-element group 507 transition  output  bypass 
    -- predecessors 488 
    -- successors 509 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_2729_to_assign_stmt_2799/AND_u32_u32_2758_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_2729_to_assign_stmt_2799/AND_u32_u32_2758_Update/cr
      -- 	branch_block_stmt_2042/assign_stmt_2729_to_assign_stmt_2799/AND_u32_u32_2758_Update/$entry
      -- 
    cp_elements(507) <= cp_elements(488);
    cr_12410_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(507), ack => AND_u32_u32_2758_inst_req_1); -- 
    -- CP-element group 508 transition  input  bypass 
    -- predecessors 506 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_2729_to_assign_stmt_2799/AND_u32_u32_2758_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2729_to_assign_stmt_2799/AND_u32_u32_2758_Sample/$exit
      -- 	branch_block_stmt_2042/assign_stmt_2729_to_assign_stmt_2799/AND_u32_u32_2758_Sample/ra
      -- 
    ra_12406_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => AND_u32_u32_2758_inst_ack_0, ack => cp_elements(508)); -- 
    -- CP-element group 509 transition  input  output  bypass 
    -- predecessors 507 
    -- successors 511 
    -- members (10) 
      -- 	branch_block_stmt_2042/assign_stmt_2729_to_assign_stmt_2799/R_iNsTr_69_2761_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_2729_to_assign_stmt_2799/R_iNsTr_69_2761_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2729_to_assign_stmt_2799/OR_u32_u32_2764_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_2729_to_assign_stmt_2799/AND_u32_u32_2758_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2729_to_assign_stmt_2799/R_iNsTr_69_2761_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2729_to_assign_stmt_2799/OR_u32_u32_2764_Sample/$entry
      -- 	branch_block_stmt_2042/assign_stmt_2729_to_assign_stmt_2799/OR_u32_u32_2764_Sample/rr
      -- 	branch_block_stmt_2042/assign_stmt_2729_to_assign_stmt_2799/AND_u32_u32_2758_Update/ca
      -- 	branch_block_stmt_2042/assign_stmt_2729_to_assign_stmt_2799/AND_u32_u32_2758_Update/$exit
      -- 	branch_block_stmt_2042/assign_stmt_2729_to_assign_stmt_2799/R_iNsTr_69_2761_update_start_
      -- 
    ca_12411_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => AND_u32_u32_2758_inst_ack_1, ack => cp_elements(509)); -- 
    rr_12423_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(509), ack => OR_u32_u32_2764_inst_req_0); -- 
    -- CP-element group 510 transition  output  bypass 
    -- predecessors 488 
    -- successors 512 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_2729_to_assign_stmt_2799/OR_u32_u32_2764_Update/$entry
      -- 	branch_block_stmt_2042/assign_stmt_2729_to_assign_stmt_2799/OR_u32_u32_2764_Update/cr
      -- 	branch_block_stmt_2042/assign_stmt_2729_to_assign_stmt_2799/OR_u32_u32_2764_update_start_
      -- 
    cp_elements(510) <= cp_elements(488);
    cr_12428_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(510), ack => OR_u32_u32_2764_inst_req_1); -- 
    -- CP-element group 511 transition  input  bypass 
    -- predecessors 509 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_2729_to_assign_stmt_2799/OR_u32_u32_2764_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2729_to_assign_stmt_2799/OR_u32_u32_2764_Sample/ra
      -- 	branch_block_stmt_2042/assign_stmt_2729_to_assign_stmt_2799/OR_u32_u32_2764_Sample/$exit
      -- 
    ra_12424_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => OR_u32_u32_2764_inst_ack_0, ack => cp_elements(511)); -- 
    -- CP-element group 512 transition  input  bypass 
    -- predecessors 510 
    -- successors 536 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_2729_to_assign_stmt_2799/OR_u32_u32_2764_Update/ca
      -- 	branch_block_stmt_2042/assign_stmt_2729_to_assign_stmt_2799/OR_u32_u32_2764_Update/$exit
      -- 	branch_block_stmt_2042/assign_stmt_2729_to_assign_stmt_2799/OR_u32_u32_2764_update_completed_
      -- 
    ca_12429_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => OR_u32_u32_2764_inst_ack_1, ack => cp_elements(512)); -- 
    -- CP-element group 513 transition  output  bypass 
    -- predecessors 488 
    -- successors 516 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_2729_to_assign_stmt_2799/LSHR_u32_u32_2770_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_2729_to_assign_stmt_2799/LSHR_u32_u32_2770_Update/$entry
      -- 	branch_block_stmt_2042/assign_stmt_2729_to_assign_stmt_2799/LSHR_u32_u32_2770_Update/cr
      -- 
    cp_elements(513) <= cp_elements(488);
    cr_12446_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(513), ack => LSHR_u32_u32_2770_inst_req_1); -- 
    -- CP-element group 514 transition  output  bypass 
    -- predecessors 488 
    -- successors 515 
    -- members (7) 
      -- 	branch_block_stmt_2042/assign_stmt_2729_to_assign_stmt_2799/LSHR_u32_u32_2770_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_2729_to_assign_stmt_2799/R_tmp6x_xix_xi2_2767_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_2729_to_assign_stmt_2799/R_tmp6x_xix_xi2_2767_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2729_to_assign_stmt_2799/R_tmp6x_xix_xi2_2767_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_2729_to_assign_stmt_2799/R_tmp6x_xix_xi2_2767_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2729_to_assign_stmt_2799/LSHR_u32_u32_2770_Sample/$entry
      -- 	branch_block_stmt_2042/assign_stmt_2729_to_assign_stmt_2799/LSHR_u32_u32_2770_Sample/rr
      -- 
    cp_elements(514) <= cp_elements(488);
    rr_12441_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(514), ack => LSHR_u32_u32_2770_inst_req_0); -- 
    -- CP-element group 515 transition  input  bypass 
    -- predecessors 514 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_2729_to_assign_stmt_2799/LSHR_u32_u32_2770_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2729_to_assign_stmt_2799/LSHR_u32_u32_2770_Sample/$exit
      -- 	branch_block_stmt_2042/assign_stmt_2729_to_assign_stmt_2799/LSHR_u32_u32_2770_Sample/ra
      -- 
    ra_12442_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => LSHR_u32_u32_2770_inst_ack_0, ack => cp_elements(515)); -- 
    -- CP-element group 516 transition  input  output  bypass 
    -- predecessors 513 
    -- successors 518 
    -- members (10) 
      -- 	branch_block_stmt_2042/assign_stmt_2729_to_assign_stmt_2799/LSHR_u32_u32_2770_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2729_to_assign_stmt_2799/LSHR_u32_u32_2770_Update/$exit
      -- 	branch_block_stmt_2042/assign_stmt_2729_to_assign_stmt_2799/LSHR_u32_u32_2770_Update/ca
      -- 	branch_block_stmt_2042/assign_stmt_2729_to_assign_stmt_2799/AND_u32_u32_2776_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_2729_to_assign_stmt_2799/R_iNsTr_71_2773_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_2729_to_assign_stmt_2799/R_iNsTr_71_2773_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2729_to_assign_stmt_2799/R_iNsTr_71_2773_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_2729_to_assign_stmt_2799/R_iNsTr_71_2773_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2729_to_assign_stmt_2799/AND_u32_u32_2776_Sample/$entry
      -- 	branch_block_stmt_2042/assign_stmt_2729_to_assign_stmt_2799/AND_u32_u32_2776_Sample/rr
      -- 
    ca_12447_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => LSHR_u32_u32_2770_inst_ack_1, ack => cp_elements(516)); -- 
    rr_12459_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(516), ack => AND_u32_u32_2776_inst_req_0); -- 
    -- CP-element group 517 transition  output  bypass 
    -- predecessors 488 
    -- successors 519 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_2729_to_assign_stmt_2799/AND_u32_u32_2776_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_2729_to_assign_stmt_2799/AND_u32_u32_2776_Update/$entry
      -- 	branch_block_stmt_2042/assign_stmt_2729_to_assign_stmt_2799/AND_u32_u32_2776_Update/cr
      -- 
    cp_elements(517) <= cp_elements(488);
    cr_12464_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(517), ack => AND_u32_u32_2776_inst_req_1); -- 
    -- CP-element group 518 transition  input  bypass 
    -- predecessors 516 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_2729_to_assign_stmt_2799/AND_u32_u32_2776_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2729_to_assign_stmt_2799/AND_u32_u32_2776_Sample/$exit
      -- 	branch_block_stmt_2042/assign_stmt_2729_to_assign_stmt_2799/AND_u32_u32_2776_Sample/ra
      -- 
    ra_12460_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => AND_u32_u32_2776_inst_ack_0, ack => cp_elements(518)); -- 
    -- CP-element group 519 transition  input  output  bypass 
    -- predecessors 517 
    -- successors 521 
    -- members (10) 
      -- 	branch_block_stmt_2042/assign_stmt_2729_to_assign_stmt_2799/AND_u32_u32_2776_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2729_to_assign_stmt_2799/AND_u32_u32_2776_Update/$exit
      -- 	branch_block_stmt_2042/assign_stmt_2729_to_assign_stmt_2799/AND_u32_u32_2776_Update/ca
      -- 	branch_block_stmt_2042/assign_stmt_2729_to_assign_stmt_2799/OR_u32_u32_2782_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_2729_to_assign_stmt_2799/R_iNsTr_72_2779_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_2729_to_assign_stmt_2799/R_iNsTr_72_2779_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2729_to_assign_stmt_2799/R_iNsTr_72_2779_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_2729_to_assign_stmt_2799/R_iNsTr_72_2779_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2729_to_assign_stmt_2799/OR_u32_u32_2782_Sample/$entry
      -- 	branch_block_stmt_2042/assign_stmt_2729_to_assign_stmt_2799/OR_u32_u32_2782_Sample/rr
      -- 
    ca_12465_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => AND_u32_u32_2776_inst_ack_1, ack => cp_elements(519)); -- 
    rr_12477_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(519), ack => OR_u32_u32_2782_inst_req_0); -- 
    -- CP-element group 520 transition  output  bypass 
    -- predecessors 488 
    -- successors 522 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_2729_to_assign_stmt_2799/OR_u32_u32_2782_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_2729_to_assign_stmt_2799/OR_u32_u32_2782_Update/$entry
      -- 	branch_block_stmt_2042/assign_stmt_2729_to_assign_stmt_2799/OR_u32_u32_2782_Update/cr
      -- 
    cp_elements(520) <= cp_elements(488);
    cr_12482_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(520), ack => OR_u32_u32_2782_inst_req_1); -- 
    -- CP-element group 521 transition  input  bypass 
    -- predecessors 519 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_2729_to_assign_stmt_2799/OR_u32_u32_2782_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2729_to_assign_stmt_2799/OR_u32_u32_2782_Sample/$exit
      -- 	branch_block_stmt_2042/assign_stmt_2729_to_assign_stmt_2799/OR_u32_u32_2782_Sample/ra
      -- 
    ra_12478_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => OR_u32_u32_2782_inst_ack_0, ack => cp_elements(521)); -- 
    -- CP-element group 522 transition  input  bypass 
    -- predecessors 520 
    -- successors 536 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_2729_to_assign_stmt_2799/OR_u32_u32_2782_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2729_to_assign_stmt_2799/OR_u32_u32_2782_Update/$exit
      -- 	branch_block_stmt_2042/assign_stmt_2729_to_assign_stmt_2799/OR_u32_u32_2782_Update/ca
      -- 
    ca_12483_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => OR_u32_u32_2782_inst_ack_1, ack => cp_elements(522)); -- 
    -- CP-element group 523 join  transition  output  bypass 
    -- predecessors 525 526 
    -- successors 527 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_2729_to_assign_stmt_2799/XOR_u32_u32_2787_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_2729_to_assign_stmt_2799/XOR_u32_u32_2787_Sample/$entry
      -- 	branch_block_stmt_2042/assign_stmt_2729_to_assign_stmt_2799/XOR_u32_u32_2787_Sample/rr
      -- 
    cp_element_group_523: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 20) := "cp_element_group_523"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(525) & cp_elements(526);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(523), clk => clk, reset => reset); --
    end block;
    rr_12499_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(523), ack => XOR_u32_u32_2787_inst_req_0); -- 
    -- CP-element group 524 transition  output  bypass 
    -- predecessors 488 
    -- successors 528 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_2729_to_assign_stmt_2799/XOR_u32_u32_2787_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_2729_to_assign_stmt_2799/XOR_u32_u32_2787_Update/$entry
      -- 	branch_block_stmt_2042/assign_stmt_2729_to_assign_stmt_2799/XOR_u32_u32_2787_Update/cr
      -- 
    cp_elements(524) <= cp_elements(488);
    cr_12504_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(524), ack => XOR_u32_u32_2787_inst_req_1); -- 
    -- CP-element group 525 transition  bypass 
    -- predecessors 488 
    -- successors 523 
    -- members (4) 
      -- 	branch_block_stmt_2042/assign_stmt_2729_to_assign_stmt_2799/R_tmp6x_xix_xi2_2785_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_2729_to_assign_stmt_2799/R_tmp6x_xix_xi2_2785_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2729_to_assign_stmt_2799/R_tmp6x_xix_xi2_2785_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_2729_to_assign_stmt_2799/R_tmp6x_xix_xi2_2785_update_completed_
      -- 
    cp_elements(525) <= cp_elements(488);
    -- CP-element group 526 transition  bypass 
    -- predecessors 488 
    -- successors 523 
    -- members (4) 
      -- 	branch_block_stmt_2042/assign_stmt_2729_to_assign_stmt_2799/R_tmp10x_xix_xi1_2786_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_2729_to_assign_stmt_2799/R_tmp10x_xix_xi1_2786_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2729_to_assign_stmt_2799/R_tmp10x_xix_xi1_2786_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_2729_to_assign_stmt_2799/R_tmp10x_xix_xi1_2786_update_completed_
      -- 
    cp_elements(526) <= cp_elements(488);
    -- CP-element group 527 transition  input  bypass 
    -- predecessors 523 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_2729_to_assign_stmt_2799/XOR_u32_u32_2787_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2729_to_assign_stmt_2799/XOR_u32_u32_2787_Sample/$exit
      -- 	branch_block_stmt_2042/assign_stmt_2729_to_assign_stmt_2799/XOR_u32_u32_2787_Sample/ra
      -- 
    ra_12500_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => XOR_u32_u32_2787_inst_ack_0, ack => cp_elements(527)); -- 
    -- CP-element group 528 transition  input  output  bypass 
    -- predecessors 524 
    -- successors 530 
    -- members (10) 
      -- 	branch_block_stmt_2042/assign_stmt_2729_to_assign_stmt_2799/XOR_u32_u32_2787_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2729_to_assign_stmt_2799/XOR_u32_u32_2787_Update/$exit
      -- 	branch_block_stmt_2042/assign_stmt_2729_to_assign_stmt_2799/XOR_u32_u32_2787_Update/ca
      -- 	branch_block_stmt_2042/assign_stmt_2729_to_assign_stmt_2799/AND_u32_u32_2793_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_2729_to_assign_stmt_2799/R_iNsTr_74_2790_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_2729_to_assign_stmt_2799/R_iNsTr_74_2790_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2729_to_assign_stmt_2799/R_iNsTr_74_2790_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_2729_to_assign_stmt_2799/R_iNsTr_74_2790_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2729_to_assign_stmt_2799/AND_u32_u32_2793_Sample/$entry
      -- 	branch_block_stmt_2042/assign_stmt_2729_to_assign_stmt_2799/AND_u32_u32_2793_Sample/rr
      -- 
    ca_12505_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => XOR_u32_u32_2787_inst_ack_1, ack => cp_elements(528)); -- 
    rr_12517_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(528), ack => AND_u32_u32_2793_inst_req_0); -- 
    -- CP-element group 529 transition  output  bypass 
    -- predecessors 488 
    -- successors 531 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_2729_to_assign_stmt_2799/AND_u32_u32_2793_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_2729_to_assign_stmt_2799/AND_u32_u32_2793_Update/$entry
      -- 	branch_block_stmt_2042/assign_stmt_2729_to_assign_stmt_2799/AND_u32_u32_2793_Update/cr
      -- 
    cp_elements(529) <= cp_elements(488);
    cr_12522_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(529), ack => AND_u32_u32_2793_inst_req_1); -- 
    -- CP-element group 530 transition  input  bypass 
    -- predecessors 528 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_2729_to_assign_stmt_2799/AND_u32_u32_2793_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2729_to_assign_stmt_2799/AND_u32_u32_2793_Sample/$exit
      -- 	branch_block_stmt_2042/assign_stmt_2729_to_assign_stmt_2799/AND_u32_u32_2793_Sample/ra
      -- 
    ra_12518_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => AND_u32_u32_2793_inst_ack_0, ack => cp_elements(530)); -- 
    -- CP-element group 531 transition  input  bypass 
    -- predecessors 529 
    -- successors 536 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_2729_to_assign_stmt_2799/AND_u32_u32_2793_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2729_to_assign_stmt_2799/AND_u32_u32_2793_Update/$exit
      -- 	branch_block_stmt_2042/assign_stmt_2729_to_assign_stmt_2799/AND_u32_u32_2793_Update/ca
      -- 
    ca_12523_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => AND_u32_u32_2793_inst_ack_1, ack => cp_elements(531)); -- 
    -- CP-element group 532 join  transition  output  bypass 
    -- predecessors 495 502 
    -- successors 534 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_2729_to_assign_stmt_2799/SUB_u32_u32_2798_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_2729_to_assign_stmt_2799/SUB_u32_u32_2798_Sample/$entry
      -- 	branch_block_stmt_2042/assign_stmt_2729_to_assign_stmt_2799/SUB_u32_u32_2798_Sample/rr
      -- 
    cp_element_group_532: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 20) := "cp_element_group_532"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(495) & cp_elements(502);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(532), clk => clk, reset => reset); --
    end block;
    rr_12539_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(532), ack => SUB_u32_u32_2798_inst_req_0); -- 
    -- CP-element group 533 transition  output  bypass 
    -- predecessors 488 
    -- successors 535 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_2729_to_assign_stmt_2799/SUB_u32_u32_2798_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_2729_to_assign_stmt_2799/SUB_u32_u32_2798_Update/$entry
      -- 	branch_block_stmt_2042/assign_stmt_2729_to_assign_stmt_2799/SUB_u32_u32_2798_Update/cr
      -- 
    cp_elements(533) <= cp_elements(488);
    cr_12544_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(533), ack => SUB_u32_u32_2798_inst_req_1); -- 
    -- CP-element group 534 transition  input  bypass 
    -- predecessors 532 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_2729_to_assign_stmt_2799/SUB_u32_u32_2798_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2729_to_assign_stmt_2799/SUB_u32_u32_2798_Sample/$exit
      -- 	branch_block_stmt_2042/assign_stmt_2729_to_assign_stmt_2799/SUB_u32_u32_2798_Sample/ra
      -- 
    ra_12540_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => SUB_u32_u32_2798_inst_ack_0, ack => cp_elements(534)); -- 
    -- CP-element group 535 transition  input  bypass 
    -- predecessors 533 
    -- successors 536 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_2729_to_assign_stmt_2799/SUB_u32_u32_2798_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2729_to_assign_stmt_2799/SUB_u32_u32_2798_Update/$exit
      -- 	branch_block_stmt_2042/assign_stmt_2729_to_assign_stmt_2799/SUB_u32_u32_2798_Update/ca
      -- 
    ca_12545_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => SUB_u32_u32_2798_inst_ack_1, ack => cp_elements(535)); -- 
    -- CP-element group 536 join  transition  bypass 
    -- predecessors 512 522 531 535 
    -- successors 28 
    -- members (1) 
      -- 	branch_block_stmt_2042/assign_stmt_2729_to_assign_stmt_2799/$exit
      -- 
    cp_element_group_536: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 20) := "cp_element_group_536"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= cp_elements(512) & cp_elements(522) & cp_elements(531) & cp_elements(535);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(536), clk => clk, reset => reset); --
    end block;
    -- CP-element group 537 transition  place  dead  bypass 
    -- predecessors 28 
    -- successors 29 
    -- members (8) 
      -- 	branch_block_stmt_2042/switch_stmt_2800__exit__
      -- 	branch_block_stmt_2042/merge_stmt_2810__entry__
      -- 	branch_block_stmt_2042/switch_stmt_2800_dead_link/$entry
      -- 	branch_block_stmt_2042/switch_stmt_2800_dead_link/$exit
      -- 	branch_block_stmt_2042/switch_stmt_2800_dead_link/dead_transition
      -- 	branch_block_stmt_2042/merge_stmt_2810_dead_link/dead_transition
      -- 	branch_block_stmt_2042/merge_stmt_2810_dead_link/$exit
      -- 	branch_block_stmt_2042/merge_stmt_2810_dead_link/$entry
      -- 
    cp_elements(537) <= false;
    -- CP-element group 538 place  bypass 
    -- predecessors 28 
    -- successors 539 
    -- members (1) 
      -- 	branch_block_stmt_2042/switch_stmt_2800__condition_check_place__
      -- 
    cp_elements(538) <= cp_elements(28);
    -- CP-element group 539 fork  transition  bypass 
    -- predecessors 538 
    -- successors 540 546 
    -- members (1) 
      -- 	branch_block_stmt_2042/switch_stmt_2800__condition_check__/$entry
      -- 
    cp_elements(539) <= cp_elements(538);
    -- CP-element group 540 fork  transition  bypass 
    -- predecessors 539 
    -- successors 541 543 
    -- members (2) 
      -- 	branch_block_stmt_2042/switch_stmt_2800__condition_check__/condition_0/$entry
      -- 	branch_block_stmt_2042/switch_stmt_2800__condition_check__/condition_0/SplitProtocol/$entry
      -- 
    cp_elements(540) <= cp_elements(539);
    -- CP-element group 541 transition  output  bypass 
    -- predecessors 540 
    -- successors 542 
    -- members (2) 
      -- 	branch_block_stmt_2042/switch_stmt_2800__condition_check__/condition_0/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_2042/switch_stmt_2800__condition_check__/condition_0/SplitProtocol/Sample/rr
      -- 
    cp_elements(541) <= cp_elements(540);
    rr_12563_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(541), ack => switch_stmt_2800_select_expr_0_req_0); -- 
    -- CP-element group 542 transition  input  bypass 
    -- predecessors 541 
    -- successors 545 
    -- members (2) 
      -- 	branch_block_stmt_2042/switch_stmt_2800__condition_check__/condition_0/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_2042/switch_stmt_2800__condition_check__/condition_0/SplitProtocol/Sample/ra
      -- 
    ra_12564_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => switch_stmt_2800_select_expr_0_ack_0, ack => cp_elements(542)); -- 
    -- CP-element group 543 transition  output  bypass 
    -- predecessors 540 
    -- successors 544 
    -- members (2) 
      -- 	branch_block_stmt_2042/switch_stmt_2800__condition_check__/condition_0/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_2042/switch_stmt_2800__condition_check__/condition_0/SplitProtocol/Update/cr
      -- 
    cp_elements(543) <= cp_elements(540);
    cr_12568_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(543), ack => switch_stmt_2800_select_expr_0_req_1); -- 
    -- CP-element group 544 transition  input  bypass 
    -- predecessors 543 
    -- successors 545 
    -- members (2) 
      -- 	branch_block_stmt_2042/switch_stmt_2800__condition_check__/condition_0/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_2042/switch_stmt_2800__condition_check__/condition_0/SplitProtocol/Update/ca
      -- 
    ca_12569_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => switch_stmt_2800_select_expr_0_ack_1, ack => cp_elements(544)); -- 
    -- CP-element group 545 join  transition  output  bypass 
    -- predecessors 542 544 
    -- successors 552 
    -- members (3) 
      -- 	branch_block_stmt_2042/switch_stmt_2800__condition_check__/condition_0/$exit
      -- 	branch_block_stmt_2042/switch_stmt_2800__condition_check__/condition_0/SplitProtocol/$exit
      -- 	branch_block_stmt_2042/switch_stmt_2800__condition_check__/condition_0/cmp
      -- 
    cp_element_group_545: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 20) := "cp_element_group_545"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(542) & cp_elements(544);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(545), clk => clk, reset => reset); --
    end block;
    cmp_12570_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(545), ack => switch_stmt_2800_branch_0_req_0); -- 
    -- CP-element group 546 fork  transition  bypass 
    -- predecessors 539 
    -- successors 547 549 
    -- members (2) 
      -- 	branch_block_stmt_2042/switch_stmt_2800__condition_check__/condition_1/$entry
      -- 	branch_block_stmt_2042/switch_stmt_2800__condition_check__/condition_1/SplitProtocol/$entry
      -- 
    cp_elements(546) <= cp_elements(539);
    -- CP-element group 547 transition  output  bypass 
    -- predecessors 546 
    -- successors 548 
    -- members (2) 
      -- 	branch_block_stmt_2042/switch_stmt_2800__condition_check__/condition_1/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_2042/switch_stmt_2800__condition_check__/condition_1/SplitProtocol/Sample/rr
      -- 
    cp_elements(547) <= cp_elements(546);
    rr_12580_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(547), ack => switch_stmt_2800_select_expr_1_req_0); -- 
    -- CP-element group 548 transition  input  bypass 
    -- predecessors 547 
    -- successors 551 
    -- members (2) 
      -- 	branch_block_stmt_2042/switch_stmt_2800__condition_check__/condition_1/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_2042/switch_stmt_2800__condition_check__/condition_1/SplitProtocol/Sample/ra
      -- 
    ra_12581_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => switch_stmt_2800_select_expr_1_ack_0, ack => cp_elements(548)); -- 
    -- CP-element group 549 transition  output  bypass 
    -- predecessors 546 
    -- successors 550 
    -- members (2) 
      -- 	branch_block_stmt_2042/switch_stmt_2800__condition_check__/condition_1/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_2042/switch_stmt_2800__condition_check__/condition_1/SplitProtocol/Update/cr
      -- 
    cp_elements(549) <= cp_elements(546);
    cr_12585_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(549), ack => switch_stmt_2800_select_expr_1_req_1); -- 
    -- CP-element group 550 transition  input  bypass 
    -- predecessors 549 
    -- successors 551 
    -- members (2) 
      -- 	branch_block_stmt_2042/switch_stmt_2800__condition_check__/condition_1/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_2042/switch_stmt_2800__condition_check__/condition_1/SplitProtocol/Update/ca
      -- 
    ca_12586_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => switch_stmt_2800_select_expr_1_ack_1, ack => cp_elements(550)); -- 
    -- CP-element group 551 join  transition  output  bypass 
    -- predecessors 548 550 
    -- successors 552 
    -- members (3) 
      -- 	branch_block_stmt_2042/switch_stmt_2800__condition_check__/condition_1/$exit
      -- 	branch_block_stmt_2042/switch_stmt_2800__condition_check__/condition_1/SplitProtocol/$exit
      -- 	branch_block_stmt_2042/switch_stmt_2800__condition_check__/condition_1/cmp
      -- 
    cp_element_group_551: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 20) := "cp_element_group_551"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(548) & cp_elements(550);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(551), clk => clk, reset => reset); --
    end block;
    cmp_12587_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(551), ack => switch_stmt_2800_branch_1_req_0); -- 
    -- CP-element group 552 join  transition  output  bypass 
    -- predecessors 545 551 
    -- successors 553 
    -- members (1) 
      -- 	branch_block_stmt_2042/switch_stmt_2800__condition_check__/$exit
      -- 
    cp_element_group_552: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 20) := "cp_element_group_552"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(545) & cp_elements(551);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(552), clk => clk, reset => reset); --
    end block;
    Xexit_12553_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(552), ack => switch_stmt_2800_branch_default_req_0); -- 
    -- CP-element group 553 branch  place  bypass 
    -- predecessors 552 
    -- successors 554 556 558 
    -- members (1) 
      -- 	branch_block_stmt_2042/switch_stmt_2800__select__
      -- 
    cp_elements(553) <= cp_elements(552);
    -- CP-element group 554 transition  bypass 
    -- predecessors 553 
    -- successors 555 
    -- members (1) 
      -- 	branch_block_stmt_2042/switch_stmt_2800_choice_0/$entry
      -- 
    cp_elements(554) <= cp_elements(553);
    -- CP-element group 555 fork  transition  place  input  bypass 
    -- predecessors 554 
    -- successors 1816 1817 
    -- members (8) 
      -- 	branch_block_stmt_2042/bb_26_xx_xloopexitx_xix_xix_xi13
      -- 	branch_block_stmt_2042/switch_stmt_2800_choice_0/$exit
      -- 	branch_block_stmt_2042/switch_stmt_2800_choice_0/ack1
      -- 	branch_block_stmt_2042/bb_26_xx_xloopexitx_xix_xix_xi13_PhiReq/$entry
      -- 	branch_block_stmt_2042/bb_26_xx_xloopexitx_xix_xix_xi13_PhiReq/phi_stmt_2939/$entry
      -- 	branch_block_stmt_2042/bb_26_xx_xloopexitx_xix_xix_xi13_PhiReq/phi_stmt_2939/phi_stmt_2939_sources/$entry
      -- 	branch_block_stmt_2042/bb_26_xx_xloopexitx_xix_xix_xi13_PhiReq/phi_stmt_2939/phi_stmt_2939_sources/type_cast_2945/$entry
      -- 	branch_block_stmt_2042/bb_26_xx_xloopexitx_xix_xix_xi13_PhiReq/phi_stmt_2939/phi_stmt_2939_sources/type_cast_2945/SplitProtocol/$entry
      -- 
    ack1_12592_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => switch_stmt_2800_branch_0_ack_1, ack => cp_elements(555)); -- 
    -- CP-element group 556 transition  bypass 
    -- predecessors 553 
    -- successors 557 
    -- members (1) 
      -- 	branch_block_stmt_2042/switch_stmt_2800_choice_1/$entry
      -- 
    cp_elements(556) <= cp_elements(553);
    -- CP-element group 557 fork  transition  place  input  bypass 
    -- predecessors 556 
    -- successors 1827 1831 
    -- members (6) 
      -- 	branch_block_stmt_2042/bb_26_udiv32x_xexitx_xpreheaderx_xix_xi16
      -- 	branch_block_stmt_2042/switch_stmt_2800_choice_1/$exit
      -- 	branch_block_stmt_2042/switch_stmt_2800_choice_1/ack1
      -- 	branch_block_stmt_2042/bb_26_udiv32x_xexitx_xpreheaderx_xix_xi16_PhiReq/$entry
      -- 	branch_block_stmt_2042/bb_26_udiv32x_xexitx_xpreheaderx_xix_xi16_PhiReq/phi_stmt_2949/$entry
      -- 	branch_block_stmt_2042/bb_26_udiv32x_xexitx_xpreheaderx_xix_xi16_PhiReq/phi_stmt_2949/phi_stmt_2949_sources/$entry
      -- 
    ack1_12597_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => switch_stmt_2800_branch_1_ack_1, ack => cp_elements(557)); -- 
    -- CP-element group 558 transition  bypass 
    -- predecessors 553 
    -- successors 559 
    -- members (1) 
      -- 	branch_block_stmt_2042/switch_stmt_2800_choice_default/$entry
      -- 
    cp_elements(558) <= cp_elements(553);
    -- CP-element group 559 transition  place  input  bypass 
    -- predecessors 558 
    -- successors 29 
    -- members (9) 
      -- 	branch_block_stmt_2042/bb_26_bbx_xnph7x_xix_xix_xi5x_xpreheader
      -- 	branch_block_stmt_2042/switch_stmt_2800_choice_default/$exit
      -- 	branch_block_stmt_2042/switch_stmt_2800_choice_default/ack0
      -- 	branch_block_stmt_2042/bb_26_bbx_xnph7x_xix_xix_xi5x_xpreheader_PhiReq/$exit
      -- 	branch_block_stmt_2042/bb_26_bbx_xnph7x_xix_xix_xi5x_xpreheader_PhiReq/$entry
      -- 	branch_block_stmt_2042/merge_stmt_2810_PhiReqMerge
      -- 	branch_block_stmt_2042/merge_stmt_2810_PhiAck/dummy
      -- 	branch_block_stmt_2042/merge_stmt_2810_PhiAck/$exit
      -- 	branch_block_stmt_2042/merge_stmt_2810_PhiAck/$entry
      -- 
    ack0_12602_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => switch_stmt_2800_branch_default_ack_0, ack => cp_elements(559)); -- 
    -- CP-element group 560 fork  transition  bypass 
    -- predecessors 30 
    -- successors 561 562 566 567 
    -- members (1) 
      -- 	branch_block_stmt_2042/assign_stmt_2832_to_assign_stmt_2837/$entry
      -- 
    cp_elements(560) <= cp_elements(30);
    -- CP-element group 561 transition  output  bypass 
    -- predecessors 560 
    -- successors 564 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_2832_to_assign_stmt_2837/LSHR_u32_u32_2831_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_2832_to_assign_stmt_2837/LSHR_u32_u32_2831_Update/$entry
      -- 	branch_block_stmt_2042/assign_stmt_2832_to_assign_stmt_2837/LSHR_u32_u32_2831_Update/cr
      -- 
    cp_elements(561) <= cp_elements(560);
    cr_12623_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(561), ack => LSHR_u32_u32_2831_inst_req_1); -- 
    -- CP-element group 562 transition  output  bypass 
    -- predecessors 560 
    -- successors 563 
    -- members (7) 
      -- 	branch_block_stmt_2042/assign_stmt_2832_to_assign_stmt_2837/LSHR_u32_u32_2831_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_2832_to_assign_stmt_2837/R_xx_x016x_xix_xix_xi3_2828_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_2832_to_assign_stmt_2837/R_xx_x016x_xix_xix_xi3_2828_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2832_to_assign_stmt_2837/R_xx_x016x_xix_xix_xi3_2828_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_2832_to_assign_stmt_2837/R_xx_x016x_xix_xix_xi3_2828_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2832_to_assign_stmt_2837/LSHR_u32_u32_2831_Sample/$entry
      -- 	branch_block_stmt_2042/assign_stmt_2832_to_assign_stmt_2837/LSHR_u32_u32_2831_Sample/rr
      -- 
    cp_elements(562) <= cp_elements(560);
    rr_12618_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(562), ack => LSHR_u32_u32_2831_inst_req_0); -- 
    -- CP-element group 563 transition  input  bypass 
    -- predecessors 562 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_2832_to_assign_stmt_2837/LSHR_u32_u32_2831_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2832_to_assign_stmt_2837/LSHR_u32_u32_2831_Sample/$exit
      -- 	branch_block_stmt_2042/assign_stmt_2832_to_assign_stmt_2837/LSHR_u32_u32_2831_Sample/ra
      -- 
    ra_12619_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => LSHR_u32_u32_2831_inst_ack_0, ack => cp_elements(563)); -- 
    -- CP-element group 564 transition  input  bypass 
    -- predecessors 561 
    -- successors 565 
    -- members (7) 
      -- 	branch_block_stmt_2042/assign_stmt_2832_to_assign_stmt_2837/LSHR_u32_u32_2831_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2832_to_assign_stmt_2837/LSHR_u32_u32_2831_Update/$exit
      -- 	branch_block_stmt_2042/assign_stmt_2832_to_assign_stmt_2837/LSHR_u32_u32_2831_Update/ca
      -- 	branch_block_stmt_2042/assign_stmt_2832_to_assign_stmt_2837/R_iNsTr_125_2834_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_2832_to_assign_stmt_2837/R_iNsTr_125_2834_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2832_to_assign_stmt_2837/R_iNsTr_125_2834_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_2832_to_assign_stmt_2837/R_iNsTr_125_2834_update_completed_
      -- 
    ca_12624_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => LSHR_u32_u32_2831_inst_ack_1, ack => cp_elements(564)); -- 
    -- CP-element group 565 join  transition  output  bypass 
    -- predecessors 564 567 
    -- successors 568 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_2832_to_assign_stmt_2837/UGT_u32_u1_2836_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_2832_to_assign_stmt_2837/UGT_u32_u1_2836_Sample/$entry
      -- 	branch_block_stmt_2042/assign_stmt_2832_to_assign_stmt_2837/UGT_u32_u1_2836_Sample/rr
      -- 
    cp_element_group_565: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 20) := "cp_element_group_565"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(564) & cp_elements(567);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(565), clk => clk, reset => reset); --
    end block;
    rr_12640_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(565), ack => UGT_u32_u1_2836_inst_req_0); -- 
    -- CP-element group 566 transition  output  bypass 
    -- predecessors 560 
    -- successors 569 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_2832_to_assign_stmt_2837/UGT_u32_u1_2836_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_2832_to_assign_stmt_2837/UGT_u32_u1_2836_Update/$entry
      -- 	branch_block_stmt_2042/assign_stmt_2832_to_assign_stmt_2837/UGT_u32_u1_2836_Update/cr
      -- 
    cp_elements(566) <= cp_elements(560);
    cr_12645_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(566), ack => UGT_u32_u1_2836_inst_req_1); -- 
    -- CP-element group 567 transition  bypass 
    -- predecessors 560 
    -- successors 565 
    -- members (4) 
      -- 	branch_block_stmt_2042/assign_stmt_2832_to_assign_stmt_2837/R_iNsTr_73_2835_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_2832_to_assign_stmt_2837/R_iNsTr_73_2835_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2832_to_assign_stmt_2837/R_iNsTr_73_2835_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_2832_to_assign_stmt_2837/R_iNsTr_73_2835_update_completed_
      -- 
    cp_elements(567) <= cp_elements(560);
    -- CP-element group 568 transition  input  bypass 
    -- predecessors 565 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_2832_to_assign_stmt_2837/UGT_u32_u1_2836_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2832_to_assign_stmt_2837/UGT_u32_u1_2836_Sample/$exit
      -- 	branch_block_stmt_2042/assign_stmt_2832_to_assign_stmt_2837/UGT_u32_u1_2836_Sample/ra
      -- 
    ra_12641_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => UGT_u32_u1_2836_inst_ack_0, ack => cp_elements(568)); -- 
    -- CP-element group 569 branch  transition  place  input  bypass 
    -- predecessors 566 
    -- successors 570 571 
    -- members (6) 
      -- 	branch_block_stmt_2042/assign_stmt_2832_to_assign_stmt_2837__exit__
      -- 	branch_block_stmt_2042/if_stmt_2838__entry__
      -- 	branch_block_stmt_2042/assign_stmt_2832_to_assign_stmt_2837/$exit
      -- 	branch_block_stmt_2042/assign_stmt_2832_to_assign_stmt_2837/UGT_u32_u1_2836_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2832_to_assign_stmt_2837/UGT_u32_u1_2836_Update/$exit
      -- 	branch_block_stmt_2042/assign_stmt_2832_to_assign_stmt_2837/UGT_u32_u1_2836_Update/ca
      -- 
    ca_12646_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => UGT_u32_u1_2836_inst_ack_1, ack => cp_elements(569)); -- 
    -- CP-element group 570 transition  place  dead  bypass 
    -- predecessors 569 
    -- successors 31 
    -- members (8) 
      -- 	branch_block_stmt_2042/merge_stmt_2844__entry__
      -- 	branch_block_stmt_2042/if_stmt_2838__exit__
      -- 	branch_block_stmt_2042/if_stmt_2838_dead_link/$entry
      -- 	branch_block_stmt_2042/if_stmt_2838_dead_link/$exit
      -- 	branch_block_stmt_2042/if_stmt_2838_dead_link/dead_transition
      -- 	branch_block_stmt_2042/merge_stmt_2844_dead_link/$entry
      -- 	branch_block_stmt_2042/merge_stmt_2844_dead_link/dead_transition
      -- 	branch_block_stmt_2042/merge_stmt_2844_dead_link/$exit
      -- 
    cp_elements(570) <= false;
    -- CP-element group 571 transition  output  bypass 
    -- predecessors 569 
    -- successors 572 
    -- members (3) 
      -- 	branch_block_stmt_2042/if_stmt_2838_eval_test/$entry
      -- 	branch_block_stmt_2042/if_stmt_2838_eval_test/$exit
      -- 	branch_block_stmt_2042/if_stmt_2838_eval_test/branch_req
      -- 
    cp_elements(571) <= cp_elements(569);
    branch_req_12654_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(571), ack => if_stmt_2838_branch_req_0); -- 
    -- CP-element group 572 branch  place  bypass 
    -- predecessors 571 
    -- successors 573 575 
    -- members (1) 
      -- 	branch_block_stmt_2042/R_iNsTr_126_2839_place
      -- 
    cp_elements(572) <= cp_elements(571);
    -- CP-element group 573 transition  bypass 
    -- predecessors 572 
    -- successors 574 
    -- members (1) 
      -- 	branch_block_stmt_2042/if_stmt_2838_if_link/$entry
      -- 
    cp_elements(573) <= cp_elements(572);
    -- CP-element group 574 transition  place  input  bypass 
    -- predecessors 573 
    -- successors 31 
    -- members (9) 
      -- 	branch_block_stmt_2042/if_stmt_2838_if_link/$exit
      -- 	branch_block_stmt_2042/if_stmt_2838_if_link/if_choice_transition
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xix_xi5_bbx_xnphx_xix_xix_xi8x_xpreheader
      -- 	branch_block_stmt_2042/merge_stmt_2844_PhiAck/$exit
      -- 	branch_block_stmt_2042/merge_stmt_2844_PhiAck/$entry
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xix_xi5_bbx_xnphx_xix_xix_xi8x_xpreheader_PhiReq/$exit
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xix_xi5_bbx_xnphx_xix_xix_xi8x_xpreheader_PhiReq/$entry
      -- 	branch_block_stmt_2042/merge_stmt_2844_PhiReqMerge
      -- 	branch_block_stmt_2042/merge_stmt_2844_PhiAck/dummy
      -- 
    if_choice_transition_12659_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2838_branch_ack_1, ack => cp_elements(574)); -- 
    -- CP-element group 575 transition  bypass 
    -- predecessors 572 
    -- successors 576 
    -- members (1) 
      -- 	branch_block_stmt_2042/if_stmt_2838_else_link/$entry
      -- 
    cp_elements(575) <= cp_elements(572);
    -- CP-element group 576 transition  place  input  bypass 
    -- predecessors 575 
    -- successors 1767 
    -- members (3) 
      -- 	branch_block_stmt_2042/if_stmt_2838_else_link/$exit
      -- 	branch_block_stmt_2042/if_stmt_2838_else_link/else_choice_transition
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xix_xi5_xx_x_crit_edgex_xix_xix_xi11
      -- 
    else_choice_transition_12663_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2838_branch_ack_0, ack => cp_elements(576)); -- 
    -- CP-element group 577 fork  transition  bypass 
    -- predecessors 32 
    -- successors 578 579 582 583 587 588 
    -- members (1) 
      -- 	branch_block_stmt_2042/assign_stmt_2866_to_assign_stmt_2877/$entry
      -- 
    cp_elements(577) <= cp_elements(32);
    -- CP-element group 578 transition  output  bypass 
    -- predecessors 577 
    -- successors 581 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_2866_to_assign_stmt_2877/SHL_u32_u32_2865_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_2866_to_assign_stmt_2877/SHL_u32_u32_2865_Update/$entry
      -- 	branch_block_stmt_2042/assign_stmt_2866_to_assign_stmt_2877/SHL_u32_u32_2865_Update/cr
      -- 
    cp_elements(578) <= cp_elements(577);
    cr_12685_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(578), ack => SHL_u32_u32_2865_inst_req_1); -- 
    -- CP-element group 579 transition  output  bypass 
    -- predecessors 577 
    -- successors 580 
    -- members (7) 
      -- 	branch_block_stmt_2042/assign_stmt_2866_to_assign_stmt_2877/SHL_u32_u32_2865_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_2866_to_assign_stmt_2877/R_shifted_divisorx_x03x_xix_xix_xi6_2862_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_2866_to_assign_stmt_2877/R_shifted_divisorx_x03x_xix_xix_xi6_2862_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2866_to_assign_stmt_2877/R_shifted_divisorx_x03x_xix_xix_xi6_2862_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_2866_to_assign_stmt_2877/R_shifted_divisorx_x03x_xix_xix_xi6_2862_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2866_to_assign_stmt_2877/SHL_u32_u32_2865_Sample/$entry
      -- 	branch_block_stmt_2042/assign_stmt_2866_to_assign_stmt_2877/SHL_u32_u32_2865_Sample/rr
      -- 
    cp_elements(579) <= cp_elements(577);
    rr_12680_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(579), ack => SHL_u32_u32_2865_inst_req_0); -- 
    -- CP-element group 580 transition  input  bypass 
    -- predecessors 579 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_2866_to_assign_stmt_2877/SHL_u32_u32_2865_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2866_to_assign_stmt_2877/SHL_u32_u32_2865_Sample/$exit
      -- 	branch_block_stmt_2042/assign_stmt_2866_to_assign_stmt_2877/SHL_u32_u32_2865_Sample/ra
      -- 
    ra_12681_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => SHL_u32_u32_2865_inst_ack_0, ack => cp_elements(580)); -- 
    -- CP-element group 581 transition  input  bypass 
    -- predecessors 578 
    -- successors 586 
    -- members (7) 
      -- 	branch_block_stmt_2042/assign_stmt_2866_to_assign_stmt_2877/SHL_u32_u32_2865_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2866_to_assign_stmt_2877/SHL_u32_u32_2865_Update/$exit
      -- 	branch_block_stmt_2042/assign_stmt_2866_to_assign_stmt_2877/SHL_u32_u32_2865_Update/ca
      -- 	branch_block_stmt_2042/assign_stmt_2866_to_assign_stmt_2877/R_iNsTr_199_2874_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_2866_to_assign_stmt_2877/R_iNsTr_199_2874_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2866_to_assign_stmt_2877/R_iNsTr_199_2874_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_2866_to_assign_stmt_2877/R_iNsTr_199_2874_update_completed_
      -- 
    ca_12686_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => SHL_u32_u32_2865_inst_ack_1, ack => cp_elements(581)); -- 
    -- CP-element group 582 transition  output  bypass 
    -- predecessors 577 
    -- successors 585 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_2866_to_assign_stmt_2877/SHL_u32_u32_2871_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_2866_to_assign_stmt_2877/SHL_u32_u32_2871_Update/$entry
      -- 	branch_block_stmt_2042/assign_stmt_2866_to_assign_stmt_2877/SHL_u32_u32_2871_Update/cr
      -- 
    cp_elements(582) <= cp_elements(577);
    cr_12703_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(582), ack => SHL_u32_u32_2871_inst_req_1); -- 
    -- CP-element group 583 transition  output  bypass 
    -- predecessors 577 
    -- successors 584 
    -- members (7) 
      -- 	branch_block_stmt_2042/assign_stmt_2866_to_assign_stmt_2877/SHL_u32_u32_2871_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_2866_to_assign_stmt_2877/R_curr_quotientx_x02x_xix_xix_xi7_2868_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_2866_to_assign_stmt_2877/R_curr_quotientx_x02x_xix_xix_xi7_2868_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2866_to_assign_stmt_2877/R_curr_quotientx_x02x_xix_xix_xi7_2868_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_2866_to_assign_stmt_2877/R_curr_quotientx_x02x_xix_xix_xi7_2868_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2866_to_assign_stmt_2877/SHL_u32_u32_2871_Sample/$entry
      -- 	branch_block_stmt_2042/assign_stmt_2866_to_assign_stmt_2877/SHL_u32_u32_2871_Sample/rr
      -- 
    cp_elements(583) <= cp_elements(577);
    rr_12698_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(583), ack => SHL_u32_u32_2871_inst_req_0); -- 
    -- CP-element group 584 transition  input  bypass 
    -- predecessors 583 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_2866_to_assign_stmt_2877/SHL_u32_u32_2871_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2866_to_assign_stmt_2877/SHL_u32_u32_2871_Sample/$exit
      -- 	branch_block_stmt_2042/assign_stmt_2866_to_assign_stmt_2877/SHL_u32_u32_2871_Sample/ra
      -- 
    ra_12699_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => SHL_u32_u32_2871_inst_ack_0, ack => cp_elements(584)); -- 
    -- CP-element group 585 transition  input  bypass 
    -- predecessors 582 
    -- successors 591 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_2866_to_assign_stmt_2877/SHL_u32_u32_2871_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2866_to_assign_stmt_2877/SHL_u32_u32_2871_Update/$exit
      -- 	branch_block_stmt_2042/assign_stmt_2866_to_assign_stmt_2877/SHL_u32_u32_2871_Update/ca
      -- 
    ca_12704_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => SHL_u32_u32_2871_inst_ack_1, ack => cp_elements(585)); -- 
    -- CP-element group 586 join  transition  output  bypass 
    -- predecessors 581 588 
    -- successors 589 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_2866_to_assign_stmt_2877/ULT_u32_u1_2876_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_2866_to_assign_stmt_2877/ULT_u32_u1_2876_Sample/$entry
      -- 	branch_block_stmt_2042/assign_stmt_2866_to_assign_stmt_2877/ULT_u32_u1_2876_Sample/rr
      -- 
    cp_element_group_586: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 20) := "cp_element_group_586"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(581) & cp_elements(588);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(586), clk => clk, reset => reset); --
    end block;
    rr_12720_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(586), ack => ULT_u32_u1_2876_inst_req_0); -- 
    -- CP-element group 587 transition  output  bypass 
    -- predecessors 577 
    -- successors 590 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_2866_to_assign_stmt_2877/ULT_u32_u1_2876_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_2866_to_assign_stmt_2877/ULT_u32_u1_2876_Update/$entry
      -- 	branch_block_stmt_2042/assign_stmt_2866_to_assign_stmt_2877/ULT_u32_u1_2876_Update/cr
      -- 
    cp_elements(587) <= cp_elements(577);
    cr_12725_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(587), ack => ULT_u32_u1_2876_inst_req_1); -- 
    -- CP-element group 588 transition  bypass 
    -- predecessors 577 
    -- successors 586 
    -- members (4) 
      -- 	branch_block_stmt_2042/assign_stmt_2866_to_assign_stmt_2877/R_iNsTr_125_2875_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_2866_to_assign_stmt_2877/R_iNsTr_125_2875_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2866_to_assign_stmt_2877/R_iNsTr_125_2875_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_2866_to_assign_stmt_2877/R_iNsTr_125_2875_update_completed_
      -- 
    cp_elements(588) <= cp_elements(577);
    -- CP-element group 589 transition  input  bypass 
    -- predecessors 586 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_2866_to_assign_stmt_2877/ULT_u32_u1_2876_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2866_to_assign_stmt_2877/ULT_u32_u1_2876_Sample/$exit
      -- 	branch_block_stmt_2042/assign_stmt_2866_to_assign_stmt_2877/ULT_u32_u1_2876_Sample/ra
      -- 
    ra_12721_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ULT_u32_u1_2876_inst_ack_0, ack => cp_elements(589)); -- 
    -- CP-element group 590 transition  input  bypass 
    -- predecessors 587 
    -- successors 591 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_2866_to_assign_stmt_2877/ULT_u32_u1_2876_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2866_to_assign_stmt_2877/ULT_u32_u1_2876_Update/$exit
      -- 	branch_block_stmt_2042/assign_stmt_2866_to_assign_stmt_2877/ULT_u32_u1_2876_Update/ca
      -- 
    ca_12726_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ULT_u32_u1_2876_inst_ack_1, ack => cp_elements(590)); -- 
    -- CP-element group 591 join  transition  bypass 
    -- predecessors 585 590 
    -- successors 33 
    -- members (1) 
      -- 	branch_block_stmt_2042/assign_stmt_2866_to_assign_stmt_2877/$exit
      -- 
    cp_element_group_591: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 20) := "cp_element_group_591"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(585) & cp_elements(590);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(591), clk => clk, reset => reset); --
    end block;
    -- CP-element group 592 transition  place  dead  bypass 
    -- predecessors 33 
    -- successors 34 
    -- members (8) 
      -- 	branch_block_stmt_2042/merge_stmt_2884__entry__
      -- 	branch_block_stmt_2042/if_stmt_2878__exit__
      -- 	branch_block_stmt_2042/if_stmt_2878_dead_link/$entry
      -- 	branch_block_stmt_2042/if_stmt_2878_dead_link/$exit
      -- 	branch_block_stmt_2042/if_stmt_2878_dead_link/dead_transition
      -- 	branch_block_stmt_2042/merge_stmt_2884_dead_link/$entry
      -- 	branch_block_stmt_2042/merge_stmt_2884_dead_link/$exit
      -- 	branch_block_stmt_2042/merge_stmt_2884_dead_link/dead_transition
      -- 
    cp_elements(592) <= false;
    -- CP-element group 593 transition  output  bypass 
    -- predecessors 33 
    -- successors 594 
    -- members (3) 
      -- 	branch_block_stmt_2042/if_stmt_2878_eval_test/$entry
      -- 	branch_block_stmt_2042/if_stmt_2878_eval_test/$exit
      -- 	branch_block_stmt_2042/if_stmt_2878_eval_test/branch_req
      -- 
    cp_elements(593) <= cp_elements(33);
    branch_req_12734_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(593), ack => if_stmt_2878_branch_req_0); -- 
    -- CP-element group 594 branch  place  bypass 
    -- predecessors 593 
    -- successors 595 597 
    -- members (1) 
      -- 	branch_block_stmt_2042/R_iNsTr_201_2879_place
      -- 
    cp_elements(594) <= cp_elements(593);
    -- CP-element group 595 transition  bypass 
    -- predecessors 594 
    -- successors 596 
    -- members (1) 
      -- 	branch_block_stmt_2042/if_stmt_2878_if_link/$entry
      -- 
    cp_elements(595) <= cp_elements(594);
    -- CP-element group 596 transition  place  input  bypass 
    -- predecessors 595 
    -- successors 1705 
    -- members (3) 
      -- 	branch_block_stmt_2042/if_stmt_2878_if_link/$exit
      -- 	branch_block_stmt_2042/if_stmt_2878_if_link/if_choice_transition
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi8_bbx_xnphx_xix_xix_xi8
      -- 
    if_choice_transition_12739_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2878_branch_ack_1, ack => cp_elements(596)); -- 
    -- CP-element group 597 transition  bypass 
    -- predecessors 594 
    -- successors 598 
    -- members (1) 
      -- 	branch_block_stmt_2042/if_stmt_2878_else_link/$entry
      -- 
    cp_elements(597) <= cp_elements(594);
    -- CP-element group 598 transition  place  input  bypass 
    -- predecessors 597 
    -- successors 1748 
    -- members (3) 
      -- 	branch_block_stmt_2042/if_stmt_2878_else_link/$exit
      -- 	branch_block_stmt_2042/if_stmt_2878_else_link/else_choice_transition
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi8_xx_x_crit_edgex_xix_xix_xi11x_xloopexit
      -- 
    else_choice_transition_12743_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2878_branch_ack_0, ack => cp_elements(598)); -- 
    -- CP-element group 599 fork  transition  bypass 
    -- predecessors 35 
    -- successors 601 602 603 607 608 609 613 614 
    -- members (1) 
      -- 	branch_block_stmt_2042/assign_stmt_2914_to_assign_stmt_2924/$entry
      -- 
    cp_elements(599) <= cp_elements(35);
    -- CP-element group 600 join  transition  output  bypass 
    -- predecessors 602 603 
    -- successors 604 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_2914_to_assign_stmt_2924/ADD_u32_u32_2913_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_2914_to_assign_stmt_2924/ADD_u32_u32_2913_Sample/$entry
      -- 	branch_block_stmt_2042/assign_stmt_2914_to_assign_stmt_2924/ADD_u32_u32_2913_Sample/rr
      -- 
    cp_element_group_600: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 20) := "cp_element_group_600"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(602) & cp_elements(603);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(600), clk => clk, reset => reset); --
    end block;
    rr_12764_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(600), ack => ADD_u32_u32_2913_inst_req_0); -- 
    -- CP-element group 601 transition  output  bypass 
    -- predecessors 599 
    -- successors 605 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_2914_to_assign_stmt_2924/ADD_u32_u32_2913_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_2914_to_assign_stmt_2924/ADD_u32_u32_2913_Update/$entry
      -- 	branch_block_stmt_2042/assign_stmt_2914_to_assign_stmt_2924/ADD_u32_u32_2913_Update/cr
      -- 
    cp_elements(601) <= cp_elements(599);
    cr_12769_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(601), ack => ADD_u32_u32_2913_inst_req_1); -- 
    -- CP-element group 602 transition  bypass 
    -- predecessors 599 
    -- successors 600 
    -- members (4) 
      -- 	branch_block_stmt_2042/assign_stmt_2914_to_assign_stmt_2924/R_curr_quotientx_x0x_xlcssax_xix_xix_xi10_2911_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_2914_to_assign_stmt_2924/R_curr_quotientx_x0x_xlcssax_xix_xix_xi10_2911_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2914_to_assign_stmt_2924/R_curr_quotientx_x0x_xlcssax_xix_xix_xi10_2911_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_2914_to_assign_stmt_2924/R_curr_quotientx_x0x_xlcssax_xix_xix_xi10_2911_update_completed_
      -- 
    cp_elements(602) <= cp_elements(599);
    -- CP-element group 603 transition  bypass 
    -- predecessors 599 
    -- successors 600 
    -- members (4) 
      -- 	branch_block_stmt_2042/assign_stmt_2914_to_assign_stmt_2924/R_quotientx_x05x_xix_xix_xi4_2912_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_2914_to_assign_stmt_2924/R_quotientx_x05x_xix_xix_xi4_2912_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2914_to_assign_stmt_2924/R_quotientx_x05x_xix_xix_xi4_2912_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_2914_to_assign_stmt_2924/R_quotientx_x05x_xix_xix_xi4_2912_update_completed_
      -- 
    cp_elements(603) <= cp_elements(599);
    -- CP-element group 604 transition  input  bypass 
    -- predecessors 600 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_2914_to_assign_stmt_2924/ADD_u32_u32_2913_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2914_to_assign_stmt_2924/ADD_u32_u32_2913_Sample/$exit
      -- 	branch_block_stmt_2042/assign_stmt_2914_to_assign_stmt_2924/ADD_u32_u32_2913_Sample/ra
      -- 
    ra_12765_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u32_u32_2913_inst_ack_0, ack => cp_elements(604)); -- 
    -- CP-element group 605 transition  input  bypass 
    -- predecessors 601 
    -- successors 617 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_2914_to_assign_stmt_2924/ADD_u32_u32_2913_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2914_to_assign_stmt_2924/ADD_u32_u32_2913_Update/$exit
      -- 	branch_block_stmt_2042/assign_stmt_2914_to_assign_stmt_2924/ADD_u32_u32_2913_Update/ca
      -- 
    ca_12770_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u32_u32_2913_inst_ack_1, ack => cp_elements(605)); -- 
    -- CP-element group 606 join  transition  output  bypass 
    -- predecessors 608 609 
    -- successors 610 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_2914_to_assign_stmt_2924/SUB_u32_u32_2918_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_2914_to_assign_stmt_2924/SUB_u32_u32_2918_Sample/$entry
      -- 	branch_block_stmt_2042/assign_stmt_2914_to_assign_stmt_2924/SUB_u32_u32_2918_Sample/rr
      -- 
    cp_element_group_606: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 20) := "cp_element_group_606"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(608) & cp_elements(609);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(606), clk => clk, reset => reset); --
    end block;
    rr_12786_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(606), ack => SUB_u32_u32_2918_inst_req_0); -- 
    -- CP-element group 607 transition  output  bypass 
    -- predecessors 599 
    -- successors 611 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_2914_to_assign_stmt_2924/SUB_u32_u32_2918_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_2914_to_assign_stmt_2924/SUB_u32_u32_2918_Update/$entry
      -- 	branch_block_stmt_2042/assign_stmt_2914_to_assign_stmt_2924/SUB_u32_u32_2918_Update/cr
      -- 
    cp_elements(607) <= cp_elements(599);
    cr_12791_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(607), ack => SUB_u32_u32_2918_inst_req_1); -- 
    -- CP-element group 608 transition  bypass 
    -- predecessors 599 
    -- successors 606 
    -- members (4) 
      -- 	branch_block_stmt_2042/assign_stmt_2914_to_assign_stmt_2924/R_xx_x016x_xix_xix_xi3_2916_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_2914_to_assign_stmt_2924/R_xx_x016x_xix_xix_xi3_2916_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2914_to_assign_stmt_2924/R_xx_x016x_xix_xix_xi3_2916_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_2914_to_assign_stmt_2924/R_xx_x016x_xix_xix_xi3_2916_update_completed_
      -- 
    cp_elements(608) <= cp_elements(599);
    -- CP-element group 609 transition  bypass 
    -- predecessors 599 
    -- successors 606 
    -- members (4) 
      -- 	branch_block_stmt_2042/assign_stmt_2914_to_assign_stmt_2924/R_shifted_divisorx_x0x_xlcssax_xix_xix_xi9_2917_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_2914_to_assign_stmt_2924/R_shifted_divisorx_x0x_xlcssax_xix_xix_xi9_2917_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2914_to_assign_stmt_2924/R_shifted_divisorx_x0x_xlcssax_xix_xix_xi9_2917_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_2914_to_assign_stmt_2924/R_shifted_divisorx_x0x_xlcssax_xix_xix_xi9_2917_update_completed_
      -- 
    cp_elements(609) <= cp_elements(599);
    -- CP-element group 610 transition  input  bypass 
    -- predecessors 606 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_2914_to_assign_stmt_2924/SUB_u32_u32_2918_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2914_to_assign_stmt_2924/SUB_u32_u32_2918_Sample/$exit
      -- 	branch_block_stmt_2042/assign_stmt_2914_to_assign_stmt_2924/SUB_u32_u32_2918_Sample/ra
      -- 
    ra_12787_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => SUB_u32_u32_2918_inst_ack_0, ack => cp_elements(610)); -- 
    -- CP-element group 611 transition  input  bypass 
    -- predecessors 607 
    -- successors 612 
    -- members (7) 
      -- 	branch_block_stmt_2042/assign_stmt_2914_to_assign_stmt_2924/SUB_u32_u32_2918_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2914_to_assign_stmt_2924/SUB_u32_u32_2918_Update/$exit
      -- 	branch_block_stmt_2042/assign_stmt_2914_to_assign_stmt_2924/SUB_u32_u32_2918_Update/ca
      -- 	branch_block_stmt_2042/assign_stmt_2914_to_assign_stmt_2924/R_iNsTr_166_2921_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_2914_to_assign_stmt_2924/R_iNsTr_166_2921_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2914_to_assign_stmt_2924/R_iNsTr_166_2921_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_2914_to_assign_stmt_2924/R_iNsTr_166_2921_update_completed_
      -- 
    ca_12792_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => SUB_u32_u32_2918_inst_ack_1, ack => cp_elements(611)); -- 
    -- CP-element group 612 join  transition  output  bypass 
    -- predecessors 611 614 
    -- successors 615 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_2914_to_assign_stmt_2924/ULT_u32_u1_2923_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_2914_to_assign_stmt_2924/ULT_u32_u1_2923_Sample/$entry
      -- 	branch_block_stmt_2042/assign_stmt_2914_to_assign_stmt_2924/ULT_u32_u1_2923_Sample/rr
      -- 
    cp_element_group_612: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 20) := "cp_element_group_612"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(611) & cp_elements(614);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(612), clk => clk, reset => reset); --
    end block;
    rr_12808_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(612), ack => ULT_u32_u1_2923_inst_req_0); -- 
    -- CP-element group 613 transition  output  bypass 
    -- predecessors 599 
    -- successors 616 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_2914_to_assign_stmt_2924/ULT_u32_u1_2923_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_2914_to_assign_stmt_2924/ULT_u32_u1_2923_Update/$entry
      -- 	branch_block_stmt_2042/assign_stmt_2914_to_assign_stmt_2924/ULT_u32_u1_2923_Update/cr
      -- 
    cp_elements(613) <= cp_elements(599);
    cr_12813_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(613), ack => ULT_u32_u1_2923_inst_req_1); -- 
    -- CP-element group 614 transition  bypass 
    -- predecessors 599 
    -- successors 612 
    -- members (4) 
      -- 	branch_block_stmt_2042/assign_stmt_2914_to_assign_stmt_2924/R_iNsTr_73_2922_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_2914_to_assign_stmt_2924/R_iNsTr_73_2922_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2914_to_assign_stmt_2924/R_iNsTr_73_2922_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_2914_to_assign_stmt_2924/R_iNsTr_73_2922_update_completed_
      -- 
    cp_elements(614) <= cp_elements(599);
    -- CP-element group 615 transition  input  bypass 
    -- predecessors 612 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_2914_to_assign_stmt_2924/ULT_u32_u1_2923_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2914_to_assign_stmt_2924/ULT_u32_u1_2923_Sample/$exit
      -- 	branch_block_stmt_2042/assign_stmt_2914_to_assign_stmt_2924/ULT_u32_u1_2923_Sample/ra
      -- 
    ra_12809_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ULT_u32_u1_2923_inst_ack_0, ack => cp_elements(615)); -- 
    -- CP-element group 616 transition  input  bypass 
    -- predecessors 613 
    -- successors 617 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_2914_to_assign_stmt_2924/ULT_u32_u1_2923_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2914_to_assign_stmt_2924/ULT_u32_u1_2923_Update/$exit
      -- 	branch_block_stmt_2042/assign_stmt_2914_to_assign_stmt_2924/ULT_u32_u1_2923_Update/ca
      -- 
    ca_12814_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ULT_u32_u1_2923_inst_ack_1, ack => cp_elements(616)); -- 
    -- CP-element group 617 join  transition  bypass 
    -- predecessors 605 616 
    -- successors 36 
    -- members (1) 
      -- 	branch_block_stmt_2042/assign_stmt_2914_to_assign_stmt_2924/$exit
      -- 
    cp_element_group_617: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 20) := "cp_element_group_617"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(605) & cp_elements(616);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(617), clk => clk, reset => reset); --
    end block;
    -- CP-element group 618 transition  place  dead  bypass 
    -- predecessors 36 
    -- successors 37 
    -- members (8) 
      -- 	branch_block_stmt_2042/merge_stmt_2931__entry__
      -- 	branch_block_stmt_2042/if_stmt_2925__exit__
      -- 	branch_block_stmt_2042/if_stmt_2925_dead_link/$entry
      -- 	branch_block_stmt_2042/if_stmt_2925_dead_link/$exit
      -- 	branch_block_stmt_2042/if_stmt_2925_dead_link/dead_transition
      -- 	branch_block_stmt_2042/merge_stmt_2931_dead_link/$entry
      -- 	branch_block_stmt_2042/merge_stmt_2931_dead_link/$exit
      -- 	branch_block_stmt_2042/merge_stmt_2931_dead_link/dead_transition
      -- 
    cp_elements(618) <= false;
    -- CP-element group 619 transition  output  bypass 
    -- predecessors 36 
    -- successors 620 
    -- members (3) 
      -- 	branch_block_stmt_2042/if_stmt_2925_eval_test/$entry
      -- 	branch_block_stmt_2042/if_stmt_2925_eval_test/$exit
      -- 	branch_block_stmt_2042/if_stmt_2925_eval_test/branch_req
      -- 
    cp_elements(619) <= cp_elements(36);
    branch_req_12822_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(619), ack => if_stmt_2925_branch_req_0); -- 
    -- CP-element group 620 branch  place  bypass 
    -- predecessors 619 
    -- successors 621 623 
    -- members (1) 
      -- 	branch_block_stmt_2042/R_iNsTr_167_2926_place
      -- 
    cp_elements(620) <= cp_elements(619);
    -- CP-element group 621 transition  bypass 
    -- predecessors 620 
    -- successors 622 
    -- members (1) 
      -- 	branch_block_stmt_2042/if_stmt_2925_if_link/$entry
      -- 
    cp_elements(621) <= cp_elements(620);
    -- CP-element group 622 fork  transition  place  input  bypass 
    -- predecessors 621 
    -- successors 1810 1812 
    -- members (8) 
      -- 	branch_block_stmt_2042/if_stmt_2925_if_link/$exit
      -- 	branch_block_stmt_2042/if_stmt_2925_if_link/if_choice_transition
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi11_xx_xloopexitx_xix_xix_xi13x_xloopexit
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi11_xx_xloopexitx_xix_xix_xi13x_xloopexit_PhiReq/$entry
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi11_xx_xloopexitx_xix_xix_xi13x_xloopexit_PhiReq/phi_stmt_2932/$entry
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi11_xx_xloopexitx_xix_xix_xi13x_xloopexit_PhiReq/phi_stmt_2932/phi_stmt_2932_sources/$entry
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi11_xx_xloopexitx_xix_xix_xi13x_xloopexit_PhiReq/phi_stmt_2932/phi_stmt_2932_sources/type_cast_2935/$entry
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi11_xx_xloopexitx_xix_xix_xi13x_xloopexit_PhiReq/phi_stmt_2932/phi_stmt_2932_sources/type_cast_2935/SplitProtocol/$entry
      -- 
    if_choice_transition_12827_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2925_branch_ack_1, ack => cp_elements(622)); -- 
    -- CP-element group 623 transition  bypass 
    -- predecessors 620 
    -- successors 624 
    -- members (1) 
      -- 	branch_block_stmt_2042/if_stmt_2925_else_link/$entry
      -- 
    cp_elements(623) <= cp_elements(620);
    -- CP-element group 624 transition  place  input  bypass 
    -- predecessors 623 
    -- successors 1680 
    -- members (3) 
      -- 	branch_block_stmt_2042/if_stmt_2925_else_link/$exit
      -- 	branch_block_stmt_2042/if_stmt_2925_else_link/else_choice_transition
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi11_bbx_xnph7x_xix_xix_xi5
      -- 
    else_choice_transition_12831_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2925_branch_ack_0, ack => cp_elements(624)); -- 
    -- CP-element group 625 fork  transition  bypass 
    -- predecessors 1851 
    -- successors 626 627 630 633 634 640 
    -- members (1) 
      -- 	branch_block_stmt_2042/assign_stmt_2961_to_assign_stmt_2980/$entry
      -- 
    cp_elements(625) <= cp_elements(1851);
    -- CP-element group 626 transition  output  bypass 
    -- predecessors 625 
    -- successors 629 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_2961_to_assign_stmt_2980/AND_u32_u32_2960_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_2961_to_assign_stmt_2980/AND_u32_u32_2960_Update/$entry
      -- 	branch_block_stmt_2042/assign_stmt_2961_to_assign_stmt_2980/AND_u32_u32_2960_Update/cr
      -- 
    cp_elements(626) <= cp_elements(625);
    cr_12853_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(626), ack => AND_u32_u32_2960_inst_req_1); -- 
    -- CP-element group 627 transition  output  bypass 
    -- predecessors 625 
    -- successors 628 
    -- members (7) 
      -- 	branch_block_stmt_2042/assign_stmt_2961_to_assign_stmt_2980/AND_u32_u32_2960_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_2961_to_assign_stmt_2980/R_tempx_x0x_xphx_xix_xi14_2957_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_2961_to_assign_stmt_2980/R_tempx_x0x_xphx_xix_xi14_2957_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2961_to_assign_stmt_2980/R_tempx_x0x_xphx_xix_xi14_2957_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_2961_to_assign_stmt_2980/R_tempx_x0x_xphx_xix_xi14_2957_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2961_to_assign_stmt_2980/AND_u32_u32_2960_Sample/$entry
      -- 	branch_block_stmt_2042/assign_stmt_2961_to_assign_stmt_2980/AND_u32_u32_2960_Sample/rr
      -- 
    cp_elements(627) <= cp_elements(625);
    rr_12848_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(627), ack => AND_u32_u32_2960_inst_req_0); -- 
    -- CP-element group 628 transition  input  bypass 
    -- predecessors 627 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_2961_to_assign_stmt_2980/AND_u32_u32_2960_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2961_to_assign_stmt_2980/AND_u32_u32_2960_Sample/$exit
      -- 	branch_block_stmt_2042/assign_stmt_2961_to_assign_stmt_2980/AND_u32_u32_2960_Sample/ra
      -- 
    ra_12849_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => AND_u32_u32_2960_inst_ack_0, ack => cp_elements(628)); -- 
    -- CP-element group 629 transition  input  output  bypass 
    -- predecessors 626 
    -- successors 631 
    -- members (10) 
      -- 	branch_block_stmt_2042/assign_stmt_2961_to_assign_stmt_2980/AND_u32_u32_2960_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2961_to_assign_stmt_2980/AND_u32_u32_2960_Update/$exit
      -- 	branch_block_stmt_2042/assign_stmt_2961_to_assign_stmt_2980/AND_u32_u32_2960_Update/ca
      -- 	branch_block_stmt_2042/assign_stmt_2961_to_assign_stmt_2980/EQ_u32_u1_2966_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_2961_to_assign_stmt_2980/R_iNsTr_104_2963_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_2961_to_assign_stmt_2980/R_iNsTr_104_2963_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2961_to_assign_stmt_2980/R_iNsTr_104_2963_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_2961_to_assign_stmt_2980/R_iNsTr_104_2963_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2961_to_assign_stmt_2980/EQ_u32_u1_2966_Sample/$entry
      -- 	branch_block_stmt_2042/assign_stmt_2961_to_assign_stmt_2980/EQ_u32_u1_2966_Sample/rr
      -- 
    ca_12854_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => AND_u32_u32_2960_inst_ack_1, ack => cp_elements(629)); -- 
    rr_12866_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(629), ack => EQ_u32_u1_2966_inst_req_0); -- 
    -- CP-element group 630 transition  output  bypass 
    -- predecessors 625 
    -- successors 632 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_2961_to_assign_stmt_2980/EQ_u32_u1_2966_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_2961_to_assign_stmt_2980/EQ_u32_u1_2966_Update/$entry
      -- 	branch_block_stmt_2042/assign_stmt_2961_to_assign_stmt_2980/EQ_u32_u1_2966_Update/cr
      -- 
    cp_elements(630) <= cp_elements(625);
    cr_12871_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(630), ack => EQ_u32_u1_2966_inst_req_1); -- 
    -- CP-element group 631 transition  input  bypass 
    -- predecessors 629 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_2961_to_assign_stmt_2980/EQ_u32_u1_2966_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2961_to_assign_stmt_2980/EQ_u32_u1_2966_Sample/$exit
      -- 	branch_block_stmt_2042/assign_stmt_2961_to_assign_stmt_2980/EQ_u32_u1_2966_Sample/ra
      -- 
    ra_12867_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u32_u1_2966_inst_ack_0, ack => cp_elements(631)); -- 
    -- CP-element group 632 transition  input  bypass 
    -- predecessors 630 
    -- successors 639 
    -- members (7) 
      -- 	branch_block_stmt_2042/assign_stmt_2961_to_assign_stmt_2980/EQ_u32_u1_2966_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2961_to_assign_stmt_2980/EQ_u32_u1_2966_Update/$exit
      -- 	branch_block_stmt_2042/assign_stmt_2961_to_assign_stmt_2980/EQ_u32_u1_2966_Update/ca
      -- 	branch_block_stmt_2042/assign_stmt_2961_to_assign_stmt_2980/R_iNsTr_105_2977_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_2961_to_assign_stmt_2980/R_iNsTr_105_2977_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2961_to_assign_stmt_2980/R_iNsTr_105_2977_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_2961_to_assign_stmt_2980/R_iNsTr_105_2977_update_completed_
      -- 
    ca_12872_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u32_u1_2966_inst_ack_1, ack => cp_elements(632)); -- 
    -- CP-element group 633 transition  output  bypass 
    -- predecessors 625 
    -- successors 638 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_2961_to_assign_stmt_2980/NEQ_i32_u1_2974_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_2961_to_assign_stmt_2980/NEQ_i32_u1_2974_Update/$entry
      -- 	branch_block_stmt_2042/assign_stmt_2961_to_assign_stmt_2980/NEQ_i32_u1_2974_Update/cr
      -- 
    cp_elements(633) <= cp_elements(625);
    cr_12903_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(633), ack => NEQ_i32_u1_2974_inst_req_1); -- 
    -- CP-element group 634 transition  output  bypass 
    -- predecessors 625 
    -- successors 635 
    -- members (7) 
      -- 	branch_block_stmt_2042/assign_stmt_2961_to_assign_stmt_2980/type_cast_2970_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_2961_to_assign_stmt_2980/R_tempx_x0x_xphx_xix_xi14_2969_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_2961_to_assign_stmt_2980/R_tempx_x0x_xphx_xix_xi14_2969_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2961_to_assign_stmt_2980/R_tempx_x0x_xphx_xix_xi14_2969_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_2961_to_assign_stmt_2980/R_tempx_x0x_xphx_xix_xi14_2969_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2961_to_assign_stmt_2980/type_cast_2970_Sample/$entry
      -- 	branch_block_stmt_2042/assign_stmt_2961_to_assign_stmt_2980/type_cast_2970_Sample/rr
      -- 
    cp_elements(634) <= cp_elements(625);
    rr_12888_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(634), ack => type_cast_2970_inst_req_0); -- 
    -- CP-element group 635 transition  input  output  bypass 
    -- predecessors 634 
    -- successors 636 
    -- members (6) 
      -- 	branch_block_stmt_2042/assign_stmt_2961_to_assign_stmt_2980/type_cast_2970_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2961_to_assign_stmt_2980/type_cast_2970_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_2961_to_assign_stmt_2980/type_cast_2970_Sample/$exit
      -- 	branch_block_stmt_2042/assign_stmt_2961_to_assign_stmt_2980/type_cast_2970_Sample/ra
      -- 	branch_block_stmt_2042/assign_stmt_2961_to_assign_stmt_2980/type_cast_2970_Update/$entry
      -- 	branch_block_stmt_2042/assign_stmt_2961_to_assign_stmt_2980/type_cast_2970_Update/cr
      -- 
    ra_12889_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2970_inst_ack_0, ack => cp_elements(635)); -- 
    cr_12893_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(635), ack => type_cast_2970_inst_req_1); -- 
    -- CP-element group 636 transition  input  output  bypass 
    -- predecessors 635 
    -- successors 637 
    -- members (6) 
      -- 	branch_block_stmt_2042/assign_stmt_2961_to_assign_stmt_2980/NEQ_i32_u1_2974_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_2961_to_assign_stmt_2980/type_cast_2970_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2961_to_assign_stmt_2980/type_cast_2970_Update/$exit
      -- 	branch_block_stmt_2042/assign_stmt_2961_to_assign_stmt_2980/type_cast_2970_Update/ca
      -- 	branch_block_stmt_2042/assign_stmt_2961_to_assign_stmt_2980/NEQ_i32_u1_2974_Sample/$entry
      -- 	branch_block_stmt_2042/assign_stmt_2961_to_assign_stmt_2980/NEQ_i32_u1_2974_Sample/rr
      -- 
    ca_12894_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2970_inst_ack_1, ack => cp_elements(636)); -- 
    rr_12898_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(636), ack => NEQ_i32_u1_2974_inst_req_0); -- 
    -- CP-element group 637 transition  input  bypass 
    -- predecessors 636 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_2961_to_assign_stmt_2980/NEQ_i32_u1_2974_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2961_to_assign_stmt_2980/NEQ_i32_u1_2974_Sample/$exit
      -- 	branch_block_stmt_2042/assign_stmt_2961_to_assign_stmt_2980/NEQ_i32_u1_2974_Sample/ra
      -- 
    ra_12899_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => NEQ_i32_u1_2974_inst_ack_0, ack => cp_elements(637)); -- 
    -- CP-element group 638 transition  input  bypass 
    -- predecessors 633 
    -- successors 639 
    -- members (7) 
      -- 	branch_block_stmt_2042/assign_stmt_2961_to_assign_stmt_2980/NEQ_i32_u1_2974_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2961_to_assign_stmt_2980/NEQ_i32_u1_2974_Update/$exit
      -- 	branch_block_stmt_2042/assign_stmt_2961_to_assign_stmt_2980/NEQ_i32_u1_2974_Update/ca
      -- 	branch_block_stmt_2042/assign_stmt_2961_to_assign_stmt_2980/R_iNsTr_106_2978_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_2961_to_assign_stmt_2980/R_iNsTr_106_2978_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2961_to_assign_stmt_2980/R_iNsTr_106_2978_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_2961_to_assign_stmt_2980/R_iNsTr_106_2978_update_completed_
      -- 
    ca_12904_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => NEQ_i32_u1_2974_inst_ack_1, ack => cp_elements(638)); -- 
    -- CP-element group 639 join  transition  output  bypass 
    -- predecessors 632 638 
    -- successors 641 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_2961_to_assign_stmt_2980/AND_u1_u1_2979_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_2961_to_assign_stmt_2980/AND_u1_u1_2979_Sample/$entry
      -- 	branch_block_stmt_2042/assign_stmt_2961_to_assign_stmt_2980/AND_u1_u1_2979_Sample/rr
      -- 
    cp_element_group_639: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 20) := "cp_element_group_639"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(632) & cp_elements(638);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(639), clk => clk, reset => reset); --
    end block;
    rr_12920_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(639), ack => AND_u1_u1_2979_inst_req_0); -- 
    -- CP-element group 640 transition  output  bypass 
    -- predecessors 625 
    -- successors 642 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_2961_to_assign_stmt_2980/AND_u1_u1_2979_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_2961_to_assign_stmt_2980/AND_u1_u1_2979_Update/$entry
      -- 	branch_block_stmt_2042/assign_stmt_2961_to_assign_stmt_2980/AND_u1_u1_2979_Update/cr
      -- 
    cp_elements(640) <= cp_elements(625);
    cr_12925_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(640), ack => AND_u1_u1_2979_inst_req_1); -- 
    -- CP-element group 641 transition  input  bypass 
    -- predecessors 639 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_2961_to_assign_stmt_2980/AND_u1_u1_2979_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2961_to_assign_stmt_2980/AND_u1_u1_2979_Sample/$exit
      -- 	branch_block_stmt_2042/assign_stmt_2961_to_assign_stmt_2980/AND_u1_u1_2979_Sample/ra
      -- 
    ra_12921_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => AND_u1_u1_2979_inst_ack_0, ack => cp_elements(641)); -- 
    -- CP-element group 642 branch  transition  place  input  bypass 
    -- predecessors 640 
    -- successors 643 644 
    -- members (6) 
      -- 	branch_block_stmt_2042/assign_stmt_2961_to_assign_stmt_2980__exit__
      -- 	branch_block_stmt_2042/if_stmt_2981__entry__
      -- 	branch_block_stmt_2042/assign_stmt_2961_to_assign_stmt_2980/$exit
      -- 	branch_block_stmt_2042/assign_stmt_2961_to_assign_stmt_2980/AND_u1_u1_2979_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_2961_to_assign_stmt_2980/AND_u1_u1_2979_Update/$exit
      -- 	branch_block_stmt_2042/assign_stmt_2961_to_assign_stmt_2980/AND_u1_u1_2979_Update/ca
      -- 
    ca_12926_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => AND_u1_u1_2979_inst_ack_1, ack => cp_elements(642)); -- 
    -- CP-element group 643 transition  place  dead  bypass 
    -- predecessors 642 
    -- successors 38 
    -- members (8) 
      -- 	branch_block_stmt_2042/if_stmt_2981__exit__
      -- 	branch_block_stmt_2042/merge_stmt_2987__entry__
      -- 	branch_block_stmt_2042/if_stmt_2981_dead_link/$entry
      -- 	branch_block_stmt_2042/if_stmt_2981_dead_link/$exit
      -- 	branch_block_stmt_2042/if_stmt_2981_dead_link/dead_transition
      -- 	branch_block_stmt_2042/merge_stmt_2987_dead_link/$entry
      -- 	branch_block_stmt_2042/merge_stmt_2987_dead_link/$exit
      -- 	branch_block_stmt_2042/merge_stmt_2987_dead_link/dead_transition
      -- 
    cp_elements(643) <= false;
    -- CP-element group 644 transition  output  bypass 
    -- predecessors 642 
    -- successors 645 
    -- members (3) 
      -- 	branch_block_stmt_2042/if_stmt_2981_eval_test/$entry
      -- 	branch_block_stmt_2042/if_stmt_2981_eval_test/$exit
      -- 	branch_block_stmt_2042/if_stmt_2981_eval_test/branch_req
      -- 
    cp_elements(644) <= cp_elements(642);
    branch_req_12934_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(644), ack => if_stmt_2981_branch_req_0); -- 
    -- CP-element group 645 branch  place  bypass 
    -- predecessors 644 
    -- successors 646 648 
    -- members (1) 
      -- 	branch_block_stmt_2042/R_orx_xcond11x_xix_xi15_2982_place
      -- 
    cp_elements(645) <= cp_elements(644);
    -- CP-element group 646 transition  bypass 
    -- predecessors 645 
    -- successors 647 
    -- members (1) 
      -- 	branch_block_stmt_2042/if_stmt_2981_if_link/$entry
      -- 
    cp_elements(646) <= cp_elements(645);
    -- CP-element group 647 transition  place  input  bypass 
    -- predecessors 646 
    -- successors 38 
    -- members (9) 
      -- 	branch_block_stmt_2042/if_stmt_2981_if_link/$exit
      -- 	branch_block_stmt_2042/if_stmt_2981_if_link/if_choice_transition
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xpreheaderx_xix_xi16_udiv32x_xexitx_xix_xi20x_xpreheader
      -- 	branch_block_stmt_2042/merge_stmt_2987_PhiReqMerge
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xpreheaderx_xix_xi16_udiv32x_xexitx_xix_xi20x_xpreheader_PhiReq/$entry
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xpreheaderx_xix_xi16_udiv32x_xexitx_xix_xi20x_xpreheader_PhiReq/$exit
      -- 	branch_block_stmt_2042/merge_stmt_2987_PhiAck/$entry
      -- 	branch_block_stmt_2042/merge_stmt_2987_PhiAck/$exit
      -- 	branch_block_stmt_2042/merge_stmt_2987_PhiAck/dummy
      -- 
    if_choice_transition_12939_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2981_branch_ack_1, ack => cp_elements(647)); -- 
    -- CP-element group 648 transition  bypass 
    -- predecessors 645 
    -- successors 649 
    -- members (1) 
      -- 	branch_block_stmt_2042/if_stmt_2981_else_link/$entry
      -- 
    cp_elements(648) <= cp_elements(645);
    -- CP-element group 649 transition  place  input  bypass 
    -- predecessors 648 
    -- successors 1914 
    -- members (3) 
      -- 	branch_block_stmt_2042/if_stmt_2981_else_link/$exit
      -- 	branch_block_stmt_2042/if_stmt_2981_else_link/else_choice_transition
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xpreheaderx_xix_xi16_xx_xcritedgex_xix_xi28
      -- 
    else_choice_transition_12943_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2981_branch_ack_0, ack => cp_elements(649)); -- 
    -- CP-element group 650 fork  transition  bypass 
    -- predecessors 39 
    -- successors 651 652 655 659 662 669 672 673 
    -- members (1) 
      -- 	branch_block_stmt_2042/assign_stmt_3009_to_assign_stmt_3040/$entry
      -- 
    cp_elements(650) <= cp_elements(39);
    -- CP-element group 651 transition  output  bypass 
    -- predecessors 650 
    -- successors 654 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_3009_to_assign_stmt_3040/SHL_u32_u32_3008_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_3009_to_assign_stmt_3040/SHL_u32_u32_3008_Update/$entry
      -- 	branch_block_stmt_2042/assign_stmt_3009_to_assign_stmt_3040/SHL_u32_u32_3008_Update/cr
      -- 
    cp_elements(651) <= cp_elements(650);
    cr_12965_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(651), ack => SHL_u32_u32_3008_inst_req_1); -- 
    -- CP-element group 652 transition  output  bypass 
    -- predecessors 650 
    -- successors 653 
    -- members (7) 
      -- 	branch_block_stmt_2042/assign_stmt_3009_to_assign_stmt_3040/SHL_u32_u32_3008_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_3009_to_assign_stmt_3040/R_tempx_x012x_xix_xi17_3005_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_3009_to_assign_stmt_3040/R_tempx_x012x_xix_xi17_3005_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3009_to_assign_stmt_3040/R_tempx_x012x_xix_xi17_3005_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_3009_to_assign_stmt_3040/R_tempx_x012x_xix_xi17_3005_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3009_to_assign_stmt_3040/SHL_u32_u32_3008_Sample/$entry
      -- 	branch_block_stmt_2042/assign_stmt_3009_to_assign_stmt_3040/SHL_u32_u32_3008_Sample/rr
      -- 
    cp_elements(652) <= cp_elements(650);
    rr_12960_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(652), ack => SHL_u32_u32_3008_inst_req_0); -- 
    -- CP-element group 653 transition  input  bypass 
    -- predecessors 652 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_3009_to_assign_stmt_3040/SHL_u32_u32_3008_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3009_to_assign_stmt_3040/SHL_u32_u32_3008_Sample/$exit
      -- 	branch_block_stmt_2042/assign_stmt_3009_to_assign_stmt_3040/SHL_u32_u32_3008_Sample/ra
      -- 
    ra_12961_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => SHL_u32_u32_3008_inst_ack_0, ack => cp_elements(653)); -- 
    -- CP-element group 654 fork  transition  input  bypass 
    -- predecessors 651 
    -- successors 656 663 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_3009_to_assign_stmt_3040/SHL_u32_u32_3008_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3009_to_assign_stmt_3040/SHL_u32_u32_3008_Update/$exit
      -- 	branch_block_stmt_2042/assign_stmt_3009_to_assign_stmt_3040/SHL_u32_u32_3008_Update/ca
      -- 
    ca_12966_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => SHL_u32_u32_3008_inst_ack_1, ack => cp_elements(654)); -- 
    -- CP-element group 655 transition  output  bypass 
    -- predecessors 650 
    -- successors 658 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_3009_to_assign_stmt_3040/AND_u32_u32_3014_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_3009_to_assign_stmt_3040/AND_u32_u32_3014_Update/$entry
      -- 	branch_block_stmt_2042/assign_stmt_3009_to_assign_stmt_3040/AND_u32_u32_3014_Update/cr
      -- 
    cp_elements(655) <= cp_elements(650);
    cr_12983_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(655), ack => AND_u32_u32_3014_inst_req_1); -- 
    -- CP-element group 656 transition  output  bypass 
    -- predecessors 654 
    -- successors 657 
    -- members (7) 
      -- 	branch_block_stmt_2042/assign_stmt_3009_to_assign_stmt_3040/AND_u32_u32_3014_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_3009_to_assign_stmt_3040/R_iNsTr_170_3011_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_3009_to_assign_stmt_3040/R_iNsTr_170_3011_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3009_to_assign_stmt_3040/R_iNsTr_170_3011_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_3009_to_assign_stmt_3040/R_iNsTr_170_3011_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3009_to_assign_stmt_3040/AND_u32_u32_3014_Sample/$entry
      -- 	branch_block_stmt_2042/assign_stmt_3009_to_assign_stmt_3040/AND_u32_u32_3014_Sample/rr
      -- 
    cp_elements(656) <= cp_elements(654);
    rr_12978_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(656), ack => AND_u32_u32_3014_inst_req_0); -- 
    -- CP-element group 657 transition  input  bypass 
    -- predecessors 656 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_3009_to_assign_stmt_3040/AND_u32_u32_3014_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3009_to_assign_stmt_3040/AND_u32_u32_3014_Sample/$exit
      -- 	branch_block_stmt_2042/assign_stmt_3009_to_assign_stmt_3040/AND_u32_u32_3014_Sample/ra
      -- 
    ra_12979_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => AND_u32_u32_3014_inst_ack_0, ack => cp_elements(657)); -- 
    -- CP-element group 658 transition  input  output  bypass 
    -- predecessors 655 
    -- successors 660 
    -- members (10) 
      -- 	branch_block_stmt_2042/assign_stmt_3009_to_assign_stmt_3040/AND_u32_u32_3014_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3009_to_assign_stmt_3040/AND_u32_u32_3014_Update/$exit
      -- 	branch_block_stmt_2042/assign_stmt_3009_to_assign_stmt_3040/AND_u32_u32_3014_Update/ca
      -- 	branch_block_stmt_2042/assign_stmt_3009_to_assign_stmt_3040/EQ_u32_u1_3020_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_3009_to_assign_stmt_3040/R_iNsTr_171_3017_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_3009_to_assign_stmt_3040/R_iNsTr_171_3017_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3009_to_assign_stmt_3040/R_iNsTr_171_3017_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_3009_to_assign_stmt_3040/R_iNsTr_171_3017_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3009_to_assign_stmt_3040/EQ_u32_u1_3020_Sample/$entry
      -- 	branch_block_stmt_2042/assign_stmt_3009_to_assign_stmt_3040/EQ_u32_u1_3020_Sample/rr
      -- 
    ca_12984_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => AND_u32_u32_3014_inst_ack_1, ack => cp_elements(658)); -- 
    rr_12996_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(658), ack => EQ_u32_u1_3020_inst_req_0); -- 
    -- CP-element group 659 transition  output  bypass 
    -- predecessors 650 
    -- successors 661 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_3009_to_assign_stmt_3040/EQ_u32_u1_3020_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_3009_to_assign_stmt_3040/EQ_u32_u1_3020_Update/$entry
      -- 	branch_block_stmt_2042/assign_stmt_3009_to_assign_stmt_3040/EQ_u32_u1_3020_Update/cr
      -- 
    cp_elements(659) <= cp_elements(650);
    cr_13001_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(659), ack => EQ_u32_u1_3020_inst_req_1); -- 
    -- CP-element group 660 transition  input  bypass 
    -- predecessors 658 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_3009_to_assign_stmt_3040/EQ_u32_u1_3020_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3009_to_assign_stmt_3040/EQ_u32_u1_3020_Sample/$exit
      -- 	branch_block_stmt_2042/assign_stmt_3009_to_assign_stmt_3040/EQ_u32_u1_3020_Sample/ra
      -- 
    ra_12997_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u32_u1_3020_inst_ack_0, ack => cp_elements(660)); -- 
    -- CP-element group 661 transition  input  bypass 
    -- predecessors 659 
    -- successors 668 
    -- members (7) 
      -- 	branch_block_stmt_2042/assign_stmt_3009_to_assign_stmt_3040/R_iNsTr_172_3031_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3009_to_assign_stmt_3040/R_iNsTr_172_3031_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_3009_to_assign_stmt_3040/R_iNsTr_172_3031_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3009_to_assign_stmt_3040/R_iNsTr_172_3031_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_3009_to_assign_stmt_3040/EQ_u32_u1_3020_Update/ca
      -- 	branch_block_stmt_2042/assign_stmt_3009_to_assign_stmt_3040/EQ_u32_u1_3020_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3009_to_assign_stmt_3040/EQ_u32_u1_3020_Update/$exit
      -- 
    ca_13002_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u32_u1_3020_inst_ack_1, ack => cp_elements(661)); -- 
    -- CP-element group 662 transition  output  bypass 
    -- predecessors 650 
    -- successors 667 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_3009_to_assign_stmt_3040/NEQ_i32_u1_3028_Update/cr
      -- 	branch_block_stmt_2042/assign_stmt_3009_to_assign_stmt_3040/NEQ_i32_u1_3028_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_3009_to_assign_stmt_3040/NEQ_i32_u1_3028_Update/$entry
      -- 
    cp_elements(662) <= cp_elements(650);
    cr_13033_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(662), ack => NEQ_i32_u1_3028_inst_req_1); -- 
    -- CP-element group 663 transition  output  bypass 
    -- predecessors 654 
    -- successors 664 
    -- members (7) 
      -- 	branch_block_stmt_2042/assign_stmt_3009_to_assign_stmt_3040/type_cast_3024_Sample/rr
      -- 	branch_block_stmt_2042/assign_stmt_3009_to_assign_stmt_3040/type_cast_3024_Sample/$entry
      -- 	branch_block_stmt_2042/assign_stmt_3009_to_assign_stmt_3040/R_iNsTr_170_3023_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3009_to_assign_stmt_3040/R_iNsTr_170_3023_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_3009_to_assign_stmt_3040/R_iNsTr_170_3023_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3009_to_assign_stmt_3040/R_iNsTr_170_3023_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_3009_to_assign_stmt_3040/type_cast_3024_sample_start_
      -- 
    cp_elements(663) <= cp_elements(654);
    rr_13018_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(663), ack => type_cast_3024_inst_req_0); -- 
    -- CP-element group 664 transition  input  output  bypass 
    -- predecessors 663 
    -- successors 665 
    -- members (6) 
      -- 	branch_block_stmt_2042/assign_stmt_3009_to_assign_stmt_3040/type_cast_3024_Update/$entry
      -- 	branch_block_stmt_2042/assign_stmt_3009_to_assign_stmt_3040/type_cast_3024_Sample/ra
      -- 	branch_block_stmt_2042/assign_stmt_3009_to_assign_stmt_3040/type_cast_3024_Sample/$exit
      -- 	branch_block_stmt_2042/assign_stmt_3009_to_assign_stmt_3040/type_cast_3024_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_3009_to_assign_stmt_3040/type_cast_3024_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3009_to_assign_stmt_3040/type_cast_3024_Update/cr
      -- 
    ra_13019_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3024_inst_ack_0, ack => cp_elements(664)); -- 
    cr_13023_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(664), ack => type_cast_3024_inst_req_1); -- 
    -- CP-element group 665 transition  input  output  bypass 
    -- predecessors 664 
    -- successors 666 
    -- members (6) 
      -- 	branch_block_stmt_2042/assign_stmt_3009_to_assign_stmt_3040/NEQ_i32_u1_3028_Sample/$entry
      -- 	branch_block_stmt_2042/assign_stmt_3009_to_assign_stmt_3040/NEQ_i32_u1_3028_Sample/rr
      -- 	branch_block_stmt_2042/assign_stmt_3009_to_assign_stmt_3040/type_cast_3024_Update/$exit
      -- 	branch_block_stmt_2042/assign_stmt_3009_to_assign_stmt_3040/type_cast_3024_Update/ca
      -- 	branch_block_stmt_2042/assign_stmt_3009_to_assign_stmt_3040/type_cast_3024_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3009_to_assign_stmt_3040/NEQ_i32_u1_3028_sample_start_
      -- 
    ca_13024_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3024_inst_ack_1, ack => cp_elements(665)); -- 
    rr_13028_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(665), ack => NEQ_i32_u1_3028_inst_req_0); -- 
    -- CP-element group 666 transition  input  bypass 
    -- predecessors 665 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_3009_to_assign_stmt_3040/NEQ_i32_u1_3028_Sample/ra
      -- 	branch_block_stmt_2042/assign_stmt_3009_to_assign_stmt_3040/NEQ_i32_u1_3028_Sample/$exit
      -- 	branch_block_stmt_2042/assign_stmt_3009_to_assign_stmt_3040/NEQ_i32_u1_3028_sample_completed_
      -- 
    ra_13029_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => NEQ_i32_u1_3028_inst_ack_0, ack => cp_elements(666)); -- 
    -- CP-element group 667 transition  input  bypass 
    -- predecessors 662 
    -- successors 668 
    -- members (7) 
      -- 	branch_block_stmt_2042/assign_stmt_3009_to_assign_stmt_3040/NEQ_i32_u1_3028_Update/$exit
      -- 	branch_block_stmt_2042/assign_stmt_3009_to_assign_stmt_3040/NEQ_i32_u1_3028_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3009_to_assign_stmt_3040/R_iNsTr_173_3032_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3009_to_assign_stmt_3040/R_iNsTr_173_3032_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_3009_to_assign_stmt_3040/R_iNsTr_173_3032_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3009_to_assign_stmt_3040/R_iNsTr_173_3032_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_3009_to_assign_stmt_3040/NEQ_i32_u1_3028_Update/ca
      -- 
    ca_13034_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => NEQ_i32_u1_3028_inst_ack_1, ack => cp_elements(667)); -- 
    -- CP-element group 668 join  transition  output  bypass 
    -- predecessors 661 667 
    -- successors 670 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_3009_to_assign_stmt_3040/AND_u1_u1_3033_Sample/rr
      -- 	branch_block_stmt_2042/assign_stmt_3009_to_assign_stmt_3040/AND_u1_u1_3033_Sample/$entry
      -- 	branch_block_stmt_2042/assign_stmt_3009_to_assign_stmt_3040/AND_u1_u1_3033_sample_start_
      -- 
    cp_element_group_668: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 20) := "cp_element_group_668"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(661) & cp_elements(667);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(668), clk => clk, reset => reset); --
    end block;
    rr_13050_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(668), ack => AND_u1_u1_3033_inst_req_0); -- 
    -- CP-element group 669 transition  output  bypass 
    -- predecessors 650 
    -- successors 671 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_3009_to_assign_stmt_3040/AND_u1_u1_3033_Update/cr
      -- 	branch_block_stmt_2042/assign_stmt_3009_to_assign_stmt_3040/AND_u1_u1_3033_Update/$entry
      -- 	branch_block_stmt_2042/assign_stmt_3009_to_assign_stmt_3040/AND_u1_u1_3033_update_start_
      -- 
    cp_elements(669) <= cp_elements(650);
    cr_13055_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(669), ack => AND_u1_u1_3033_inst_req_1); -- 
    -- CP-element group 670 transition  input  bypass 
    -- predecessors 668 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_3009_to_assign_stmt_3040/AND_u1_u1_3033_Sample/ra
      -- 	branch_block_stmt_2042/assign_stmt_3009_to_assign_stmt_3040/AND_u1_u1_3033_Sample/$exit
      -- 	branch_block_stmt_2042/assign_stmt_3009_to_assign_stmt_3040/AND_u1_u1_3033_sample_completed_
      -- 
    ra_13051_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => AND_u1_u1_3033_inst_ack_0, ack => cp_elements(670)); -- 
    -- CP-element group 671 transition  input  bypass 
    -- predecessors 669 
    -- successors 676 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_3009_to_assign_stmt_3040/AND_u1_u1_3033_Update/ca
      -- 	branch_block_stmt_2042/assign_stmt_3009_to_assign_stmt_3040/AND_u1_u1_3033_Update/$exit
      -- 	branch_block_stmt_2042/assign_stmt_3009_to_assign_stmt_3040/AND_u1_u1_3033_update_completed_
      -- 
    ca_13056_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => AND_u1_u1_3033_inst_ack_1, ack => cp_elements(671)); -- 
    -- CP-element group 672 transition  output  bypass 
    -- predecessors 650 
    -- successors 675 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_3009_to_assign_stmt_3040/ADD_u32_u32_3039_Update/cr
      -- 	branch_block_stmt_2042/assign_stmt_3009_to_assign_stmt_3040/ADD_u32_u32_3039_Update/$entry
      -- 	branch_block_stmt_2042/assign_stmt_3009_to_assign_stmt_3040/ADD_u32_u32_3039_update_start_
      -- 
    cp_elements(672) <= cp_elements(650);
    cr_13073_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(672), ack => ADD_u32_u32_3039_inst_req_1); -- 
    -- CP-element group 673 transition  output  bypass 
    -- predecessors 650 
    -- successors 674 
    -- members (7) 
      -- 	branch_block_stmt_2042/assign_stmt_3009_to_assign_stmt_3040/ADD_u32_u32_3039_Sample/rr
      -- 	branch_block_stmt_2042/assign_stmt_3009_to_assign_stmt_3040/ADD_u32_u32_3039_Sample/$entry
      -- 	branch_block_stmt_2042/assign_stmt_3009_to_assign_stmt_3040/R_iNsTr_169_3036_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3009_to_assign_stmt_3040/R_iNsTr_169_3036_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_3009_to_assign_stmt_3040/R_iNsTr_169_3036_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3009_to_assign_stmt_3040/R_iNsTr_169_3036_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_3009_to_assign_stmt_3040/ADD_u32_u32_3039_sample_start_
      -- 
    cp_elements(673) <= cp_elements(650);
    rr_13068_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(673), ack => ADD_u32_u32_3039_inst_req_0); -- 
    -- CP-element group 674 transition  input  bypass 
    -- predecessors 673 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_3009_to_assign_stmt_3040/ADD_u32_u32_3039_Sample/ra
      -- 	branch_block_stmt_2042/assign_stmt_3009_to_assign_stmt_3040/ADD_u32_u32_3039_Sample/$exit
      -- 	branch_block_stmt_2042/assign_stmt_3009_to_assign_stmt_3040/ADD_u32_u32_3039_sample_completed_
      -- 
    ra_13069_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u32_u32_3039_inst_ack_0, ack => cp_elements(674)); -- 
    -- CP-element group 675 transition  input  bypass 
    -- predecessors 672 
    -- successors 676 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_3009_to_assign_stmt_3040/ADD_u32_u32_3039_Update/ca
      -- 	branch_block_stmt_2042/assign_stmt_3009_to_assign_stmt_3040/ADD_u32_u32_3039_Update/$exit
      -- 	branch_block_stmt_2042/assign_stmt_3009_to_assign_stmt_3040/ADD_u32_u32_3039_update_completed_
      -- 
    ca_13074_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u32_u32_3039_inst_ack_1, ack => cp_elements(675)); -- 
    -- CP-element group 676 join  transition  bypass 
    -- predecessors 671 675 
    -- successors 40 
    -- members (1) 
      -- 	branch_block_stmt_2042/assign_stmt_3009_to_assign_stmt_3040/$exit
      -- 
    cp_element_group_676: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 20) := "cp_element_group_676"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(671) & cp_elements(675);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(676), clk => clk, reset => reset); --
    end block;
    -- CP-element group 677 transition  place  dead  bypass 
    -- predecessors 40 
    -- successors 41 
    -- members (8) 
      -- 	branch_block_stmt_2042/merge_stmt_3047__entry__
      -- 	branch_block_stmt_2042/if_stmt_3041__exit__
      -- 	branch_block_stmt_2042/if_stmt_3041_dead_link/dead_transition
      -- 	branch_block_stmt_2042/if_stmt_3041_dead_link/$exit
      -- 	branch_block_stmt_2042/if_stmt_3041_dead_link/$entry
      -- 	branch_block_stmt_2042/merge_stmt_3047_dead_link/$entry
      -- 	branch_block_stmt_2042/merge_stmt_3047_dead_link/$exit
      -- 	branch_block_stmt_2042/merge_stmt_3047_dead_link/dead_transition
      -- 
    cp_elements(677) <= false;
    -- CP-element group 678 transition  output  bypass 
    -- predecessors 40 
    -- successors 679 
    -- members (3) 
      -- 	branch_block_stmt_2042/if_stmt_3041_eval_test/branch_req
      -- 	branch_block_stmt_2042/if_stmt_3041_eval_test/$exit
      -- 	branch_block_stmt_2042/if_stmt_3041_eval_test/$entry
      -- 
    cp_elements(678) <= cp_elements(40);
    branch_req_13082_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(678), ack => if_stmt_3041_branch_req_0); -- 
    -- CP-element group 679 branch  place  bypass 
    -- predecessors 678 
    -- successors 680 682 
    -- members (1) 
      -- 	branch_block_stmt_2042/R_orx_xcondx_xix_xi18_3042_place
      -- 
    cp_elements(679) <= cp_elements(678);
    -- CP-element group 680 transition  bypass 
    -- predecessors 679 
    -- successors 681 
    -- members (1) 
      -- 	branch_block_stmt_2042/if_stmt_3041_if_link/$entry
      -- 
    cp_elements(680) <= cp_elements(679);
    -- CP-element group 681 transition  place  input  bypass 
    -- predecessors 680 
    -- successors 1852 
    -- members (3) 
      -- 	branch_block_stmt_2042/if_stmt_3041_if_link/if_choice_transition
      -- 	branch_block_stmt_2042/if_stmt_3041_if_link/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi20_udiv32x_xexitx_xix_xi20
      -- 
    if_choice_transition_13087_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_3041_branch_ack_1, ack => cp_elements(681)); -- 
    -- CP-element group 682 transition  bypass 
    -- predecessors 679 
    -- successors 683 
    -- members (1) 
      -- 	branch_block_stmt_2042/if_stmt_3041_else_link/$entry
      -- 
    cp_elements(682) <= cp_elements(679);
    -- CP-element group 683 transition  place  input  bypass 
    -- predecessors 682 
    -- successors 1895 
    -- members (3) 
      -- 	branch_block_stmt_2042/if_stmt_3041_else_link/else_choice_transition
      -- 	branch_block_stmt_2042/if_stmt_3041_else_link/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi20_udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi24
      -- 
    else_choice_transition_13091_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_3041_branch_ack_0, ack => cp_elements(683)); -- 
    -- CP-element group 684 fork  transition  bypass 
    -- predecessors 41 
    -- successors 685 686 690 691 695 696 
    -- members (1) 
      -- 	branch_block_stmt_2042/assign_stmt_3062_to_assign_stmt_3072/$entry
      -- 
    cp_elements(684) <= cp_elements(41);
    -- CP-element group 685 transition  output  bypass 
    -- predecessors 684 
    -- successors 688 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_3062_to_assign_stmt_3072/ADD_u32_u32_3061_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_3062_to_assign_stmt_3072/ADD_u32_u32_3061_Update/$entry
      -- 	branch_block_stmt_2042/assign_stmt_3062_to_assign_stmt_3072/ADD_u32_u32_3061_Update/cr
      -- 
    cp_elements(685) <= cp_elements(684);
    cr_13113_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(685), ack => ADD_u32_u32_3061_inst_req_1); -- 
    -- CP-element group 686 transition  output  bypass 
    -- predecessors 684 
    -- successors 687 
    -- members (7) 
      -- 	branch_block_stmt_2042/assign_stmt_3062_to_assign_stmt_3072/R_iNsTr_65_3058_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_3062_to_assign_stmt_3072/R_iNsTr_65_3058_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3062_to_assign_stmt_3072/R_iNsTr_65_3058_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_3062_to_assign_stmt_3072/R_iNsTr_65_3058_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3062_to_assign_stmt_3072/ADD_u32_u32_3061_Sample/$entry
      -- 	branch_block_stmt_2042/assign_stmt_3062_to_assign_stmt_3072/ADD_u32_u32_3061_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_3062_to_assign_stmt_3072/ADD_u32_u32_3061_Sample/rr
      -- 
    cp_elements(686) <= cp_elements(684);
    rr_13108_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(686), ack => ADD_u32_u32_3061_inst_req_0); -- 
    -- CP-element group 687 transition  input  bypass 
    -- predecessors 686 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_3062_to_assign_stmt_3072/ADD_u32_u32_3061_Sample/ra
      -- 	branch_block_stmt_2042/assign_stmt_3062_to_assign_stmt_3072/ADD_u32_u32_3061_Sample/$exit
      -- 	branch_block_stmt_2042/assign_stmt_3062_to_assign_stmt_3072/ADD_u32_u32_3061_sample_completed_
      -- 
    ra_13109_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u32_u32_3061_inst_ack_0, ack => cp_elements(687)); -- 
    -- CP-element group 688 transition  input  bypass 
    -- predecessors 685 
    -- successors 689 
    -- members (7) 
      -- 	branch_block_stmt_2042/assign_stmt_3062_to_assign_stmt_3072/ADD_u32_u32_3061_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3062_to_assign_stmt_3072/ADD_u32_u32_3061_Update/$exit
      -- 	branch_block_stmt_2042/assign_stmt_3062_to_assign_stmt_3072/ADD_u32_u32_3061_Update/ca
      -- 	branch_block_stmt_2042/assign_stmt_3062_to_assign_stmt_3072/R_tmp21x_xix_xi21_3064_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3062_to_assign_stmt_3072/R_tmp21x_xix_xi21_3064_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_3062_to_assign_stmt_3072/R_tmp21x_xix_xi21_3064_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3062_to_assign_stmt_3072/R_tmp21x_xix_xi21_3064_sample_start_
      -- 
    ca_13114_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u32_u32_3061_inst_ack_1, ack => cp_elements(688)); -- 
    -- CP-element group 689 join  transition  output  bypass 
    -- predecessors 688 691 
    -- successors 692 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_3062_to_assign_stmt_3072/SUB_u32_u32_3066_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_3062_to_assign_stmt_3072/SUB_u32_u32_3066_Sample/$entry
      -- 	branch_block_stmt_2042/assign_stmt_3062_to_assign_stmt_3072/SUB_u32_u32_3066_Sample/rr
      -- 
    cp_element_group_689: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 20) := "cp_element_group_689"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(688) & cp_elements(691);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(689), clk => clk, reset => reset); --
    end block;
    rr_13130_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(689), ack => SUB_u32_u32_3066_inst_req_0); -- 
    -- CP-element group 690 transition  output  bypass 
    -- predecessors 684 
    -- successors 693 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_3062_to_assign_stmt_3072/SUB_u32_u32_3066_Update/cr
      -- 	branch_block_stmt_2042/assign_stmt_3062_to_assign_stmt_3072/SUB_u32_u32_3066_Update/$entry
      -- 	branch_block_stmt_2042/assign_stmt_3062_to_assign_stmt_3072/SUB_u32_u32_3066_update_start_
      -- 
    cp_elements(690) <= cp_elements(684);
    cr_13135_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(690), ack => SUB_u32_u32_3066_inst_req_1); -- 
    -- CP-element group 691 transition  bypass 
    -- predecessors 684 
    -- successors 689 
    -- members (4) 
      -- 	branch_block_stmt_2042/assign_stmt_3062_to_assign_stmt_3072/R_iNsTr_67_3065_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_3062_to_assign_stmt_3072/R_iNsTr_67_3065_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3062_to_assign_stmt_3072/R_iNsTr_67_3065_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3062_to_assign_stmt_3072/R_iNsTr_67_3065_sample_start_
      -- 
    cp_elements(691) <= cp_elements(684);
    -- CP-element group 692 transition  input  bypass 
    -- predecessors 689 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_3062_to_assign_stmt_3072/SUB_u32_u32_3066_Sample/$exit
      -- 	branch_block_stmt_2042/assign_stmt_3062_to_assign_stmt_3072/SUB_u32_u32_3066_Sample/ra
      -- 	branch_block_stmt_2042/assign_stmt_3062_to_assign_stmt_3072/SUB_u32_u32_3066_sample_completed_
      -- 
    ra_13131_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => SUB_u32_u32_3066_inst_ack_0, ack => cp_elements(692)); -- 
    -- CP-element group 693 transition  input  bypass 
    -- predecessors 690 
    -- successors 694 
    -- members (7) 
      -- 	branch_block_stmt_2042/assign_stmt_3062_to_assign_stmt_3072/R_tmp25x_xix_xi22_3069_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3062_to_assign_stmt_3072/SUB_u32_u32_3066_Update/$exit
      -- 	branch_block_stmt_2042/assign_stmt_3062_to_assign_stmt_3072/R_tmp25x_xix_xi22_3069_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_3062_to_assign_stmt_3072/R_tmp25x_xix_xi22_3069_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3062_to_assign_stmt_3072/R_tmp25x_xix_xi22_3069_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_3062_to_assign_stmt_3072/SUB_u32_u32_3066_Update/ca
      -- 	branch_block_stmt_2042/assign_stmt_3062_to_assign_stmt_3072/SUB_u32_u32_3066_update_completed_
      -- 
    ca_13136_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => SUB_u32_u32_3066_inst_ack_1, ack => cp_elements(693)); -- 
    -- CP-element group 694 join  transition  output  bypass 
    -- predecessors 693 696 
    -- successors 697 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_3062_to_assign_stmt_3072/SUB_u32_u32_3071_Sample/rr
      -- 	branch_block_stmt_2042/assign_stmt_3062_to_assign_stmt_3072/SUB_u32_u32_3071_Sample/$entry
      -- 	branch_block_stmt_2042/assign_stmt_3062_to_assign_stmt_3072/SUB_u32_u32_3071_sample_start_
      -- 
    cp_element_group_694: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 20) := "cp_element_group_694"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(693) & cp_elements(696);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(694), clk => clk, reset => reset); --
    end block;
    rr_13152_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(694), ack => SUB_u32_u32_3071_inst_req_0); -- 
    -- CP-element group 695 transition  output  bypass 
    -- predecessors 684 
    -- successors 698 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_3062_to_assign_stmt_3072/SUB_u32_u32_3071_Update/$entry
      -- 	branch_block_stmt_2042/assign_stmt_3062_to_assign_stmt_3072/SUB_u32_u32_3071_Update/cr
      -- 	branch_block_stmt_2042/assign_stmt_3062_to_assign_stmt_3072/SUB_u32_u32_3071_update_start_
      -- 
    cp_elements(695) <= cp_elements(684);
    cr_13157_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(695), ack => SUB_u32_u32_3071_inst_req_1); -- 
    -- CP-element group 696 transition  bypass 
    -- predecessors 684 
    -- successors 694 
    -- members (4) 
      -- 	branch_block_stmt_2042/assign_stmt_3062_to_assign_stmt_3072/R_xx_xlcssa10_3070_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_3062_to_assign_stmt_3072/R_xx_xlcssa10_3070_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3062_to_assign_stmt_3072/R_xx_xlcssa10_3070_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_3062_to_assign_stmt_3072/R_xx_xlcssa10_3070_sample_completed_
      -- 
    cp_elements(696) <= cp_elements(684);
    -- CP-element group 697 transition  input  bypass 
    -- predecessors 694 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_3062_to_assign_stmt_3072/SUB_u32_u32_3071_Sample/ra
      -- 	branch_block_stmt_2042/assign_stmt_3062_to_assign_stmt_3072/SUB_u32_u32_3071_Sample/$exit
      -- 	branch_block_stmt_2042/assign_stmt_3062_to_assign_stmt_3072/SUB_u32_u32_3071_sample_completed_
      -- 
    ra_13153_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => SUB_u32_u32_3071_inst_ack_0, ack => cp_elements(697)); -- 
    -- CP-element group 698 transition  place  input  bypass 
    -- predecessors 695 
    -- successors 1940 
    -- members (6) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi24_xx_xcritedgex_xix_xi28
      -- 	branch_block_stmt_2042/assign_stmt_3062_to_assign_stmt_3072__exit__
      -- 	branch_block_stmt_2042/assign_stmt_3062_to_assign_stmt_3072/$exit
      -- 	branch_block_stmt_2042/assign_stmt_3062_to_assign_stmt_3072/SUB_u32_u32_3071_Update/$exit
      -- 	branch_block_stmt_2042/assign_stmt_3062_to_assign_stmt_3072/SUB_u32_u32_3071_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3062_to_assign_stmt_3072/SUB_u32_u32_3071_Update/ca
      -- 
    ca_13158_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => SUB_u32_u32_3071_inst_ack_1, ack => cp_elements(698)); -- 
    -- CP-element group 699 fork  transition  bypass 
    -- predecessors 42 
    -- successors 700 701 704 705 708 712 713 717 720 
    -- members (1) 
      -- 	branch_block_stmt_2042/assign_stmt_3093_to_assign_stmt_3119/$entry
      -- 
    cp_elements(699) <= cp_elements(42);
    -- CP-element group 700 transition  output  bypass 
    -- predecessors 699 
    -- successors 703 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_3093_to_assign_stmt_3119/AND_u32_u32_3092_Update/cr
      -- 	branch_block_stmt_2042/assign_stmt_3093_to_assign_stmt_3119/AND_u32_u32_3092_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_3093_to_assign_stmt_3119/AND_u32_u32_3092_Update/$entry
      -- 
    cp_elements(700) <= cp_elements(699);
    cr_13178_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(700), ack => AND_u32_u32_3092_inst_req_1); -- 
    -- CP-element group 701 transition  output  bypass 
    -- predecessors 699 
    -- successors 702 
    -- members (7) 
      -- 	branch_block_stmt_2042/assign_stmt_3093_to_assign_stmt_3119/R_tempx_x0x_xlcssax_xix_xi26_3089_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_3093_to_assign_stmt_3119/R_tempx_x0x_xlcssax_xix_xi26_3089_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3093_to_assign_stmt_3119/R_tempx_x0x_xlcssax_xix_xi26_3089_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_3093_to_assign_stmt_3119/AND_u32_u32_3092_Sample/rr
      -- 	branch_block_stmt_2042/assign_stmt_3093_to_assign_stmt_3119/AND_u32_u32_3092_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_3093_to_assign_stmt_3119/AND_u32_u32_3092_Sample/$entry
      -- 	branch_block_stmt_2042/assign_stmt_3093_to_assign_stmt_3119/R_tempx_x0x_xlcssax_xix_xi26_3089_update_completed_
      -- 
    cp_elements(701) <= cp_elements(699);
    rr_13173_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(701), ack => AND_u32_u32_3092_inst_req_0); -- 
    -- CP-element group 702 transition  input  bypass 
    -- predecessors 701 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_3093_to_assign_stmt_3119/AND_u32_u32_3092_Sample/ra
      -- 	branch_block_stmt_2042/assign_stmt_3093_to_assign_stmt_3119/AND_u32_u32_3092_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3093_to_assign_stmt_3119/AND_u32_u32_3092_Sample/$exit
      -- 
    ra_13174_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => AND_u32_u32_3092_inst_ack_0, ack => cp_elements(702)); -- 
    -- CP-element group 703 transition  input  bypass 
    -- predecessors 700 
    -- successors 711 
    -- members (7) 
      -- 	branch_block_stmt_2042/assign_stmt_3093_to_assign_stmt_3119/R_iNsTr_129_3107_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3093_to_assign_stmt_3119/R_iNsTr_129_3107_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_3093_to_assign_stmt_3119/R_iNsTr_129_3107_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3093_to_assign_stmt_3119/R_iNsTr_129_3107_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_3093_to_assign_stmt_3119/AND_u32_u32_3092_Update/$exit
      -- 	branch_block_stmt_2042/assign_stmt_3093_to_assign_stmt_3119/AND_u32_u32_3092_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3093_to_assign_stmt_3119/AND_u32_u32_3092_Update/ca
      -- 
    ca_13179_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => AND_u32_u32_3092_inst_ack_1, ack => cp_elements(703)); -- 
    -- CP-element group 704 transition  output  bypass 
    -- predecessors 699 
    -- successors 707 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_3093_to_assign_stmt_3119/SHL_u32_u32_3098_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_3093_to_assign_stmt_3119/SHL_u32_u32_3098_Update/cr
      -- 	branch_block_stmt_2042/assign_stmt_3093_to_assign_stmt_3119/SHL_u32_u32_3098_Update/$entry
      -- 
    cp_elements(704) <= cp_elements(699);
    cr_13196_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(704), ack => SHL_u32_u32_3098_inst_req_1); -- 
    -- CP-element group 705 transition  output  bypass 
    -- predecessors 699 
    -- successors 706 
    -- members (7) 
      -- 	branch_block_stmt_2042/assign_stmt_3093_to_assign_stmt_3119/SHL_u32_u32_3098_Sample/$entry
      -- 	branch_block_stmt_2042/assign_stmt_3093_to_assign_stmt_3119/SHL_u32_u32_3098_Sample/rr
      -- 	branch_block_stmt_2042/assign_stmt_3093_to_assign_stmt_3119/R_expx_x0x_xlcssax_xix_xi25_3095_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3093_to_assign_stmt_3119/R_expx_x0x_xlcssax_xix_xi25_3095_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_3093_to_assign_stmt_3119/R_expx_x0x_xlcssax_xix_xi25_3095_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3093_to_assign_stmt_3119/R_expx_x0x_xlcssax_xix_xi25_3095_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_3093_to_assign_stmt_3119/SHL_u32_u32_3098_sample_start_
      -- 
    cp_elements(705) <= cp_elements(699);
    rr_13191_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(705), ack => SHL_u32_u32_3098_inst_req_0); -- 
    -- CP-element group 706 transition  input  bypass 
    -- predecessors 705 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_3093_to_assign_stmt_3119/SHL_u32_u32_3098_Sample/$exit
      -- 	branch_block_stmt_2042/assign_stmt_3093_to_assign_stmt_3119/SHL_u32_u32_3098_Sample/ra
      -- 	branch_block_stmt_2042/assign_stmt_3093_to_assign_stmt_3119/SHL_u32_u32_3098_sample_completed_
      -- 
    ra_13192_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => SHL_u32_u32_3098_inst_ack_0, ack => cp_elements(706)); -- 
    -- CP-element group 707 transition  input  output  bypass 
    -- predecessors 704 
    -- successors 709 
    -- members (10) 
      -- 	branch_block_stmt_2042/assign_stmt_3093_to_assign_stmt_3119/ADD_u32_u32_3104_Sample/rr
      -- 	branch_block_stmt_2042/assign_stmt_3093_to_assign_stmt_3119/ADD_u32_u32_3104_Sample/$entry
      -- 	branch_block_stmt_2042/assign_stmt_3093_to_assign_stmt_3119/R_iNsTr_130_3101_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3093_to_assign_stmt_3119/R_iNsTr_130_3101_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_3093_to_assign_stmt_3119/R_iNsTr_130_3101_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3093_to_assign_stmt_3119/R_iNsTr_130_3101_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_3093_to_assign_stmt_3119/SHL_u32_u32_3098_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3093_to_assign_stmt_3119/ADD_u32_u32_3104_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_3093_to_assign_stmt_3119/SHL_u32_u32_3098_Update/ca
      -- 	branch_block_stmt_2042/assign_stmt_3093_to_assign_stmt_3119/SHL_u32_u32_3098_Update/$exit
      -- 
    ca_13197_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => SHL_u32_u32_3098_inst_ack_1, ack => cp_elements(707)); -- 
    rr_13209_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(707), ack => ADD_u32_u32_3104_inst_req_0); -- 
    -- CP-element group 708 transition  output  bypass 
    -- predecessors 699 
    -- successors 710 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_3093_to_assign_stmt_3119/ADD_u32_u32_3104_Update/cr
      -- 	branch_block_stmt_2042/assign_stmt_3093_to_assign_stmt_3119/ADD_u32_u32_3104_Update/$entry
      -- 	branch_block_stmt_2042/assign_stmt_3093_to_assign_stmt_3119/ADD_u32_u32_3104_update_start_
      -- 
    cp_elements(708) <= cp_elements(699);
    cr_13214_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(708), ack => ADD_u32_u32_3104_inst_req_1); -- 
    -- CP-element group 709 transition  input  bypass 
    -- predecessors 707 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_3093_to_assign_stmt_3119/ADD_u32_u32_3104_Sample/ra
      -- 	branch_block_stmt_2042/assign_stmt_3093_to_assign_stmt_3119/ADD_u32_u32_3104_Sample/$exit
      -- 	branch_block_stmt_2042/assign_stmt_3093_to_assign_stmt_3119/ADD_u32_u32_3104_sample_completed_
      -- 
    ra_13210_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u32_u32_3104_inst_ack_0, ack => cp_elements(709)); -- 
    -- CP-element group 710 transition  input  bypass 
    -- predecessors 708 
    -- successors 716 
    -- members (7) 
      -- 	branch_block_stmt_2042/assign_stmt_3093_to_assign_stmt_3119/R_iNsTr_131_3113_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_3093_to_assign_stmt_3119/ADD_u32_u32_3104_Update/ca
      -- 	branch_block_stmt_2042/assign_stmt_3093_to_assign_stmt_3119/ADD_u32_u32_3104_Update/$exit
      -- 	branch_block_stmt_2042/assign_stmt_3093_to_assign_stmt_3119/R_iNsTr_131_3113_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3093_to_assign_stmt_3119/ADD_u32_u32_3104_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3093_to_assign_stmt_3119/R_iNsTr_131_3113_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3093_to_assign_stmt_3119/R_iNsTr_131_3113_update_start_
      -- 
    ca_13215_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u32_u32_3104_inst_ack_1, ack => cp_elements(710)); -- 
    -- CP-element group 711 join  transition  output  bypass 
    -- predecessors 703 713 
    -- successors 714 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_3093_to_assign_stmt_3119/OR_u32_u32_3109_Sample/rr
      -- 	branch_block_stmt_2042/assign_stmt_3093_to_assign_stmt_3119/OR_u32_u32_3109_Sample/$entry
      -- 	branch_block_stmt_2042/assign_stmt_3093_to_assign_stmt_3119/OR_u32_u32_3109_sample_start_
      -- 
    cp_element_group_711: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 20) := "cp_element_group_711"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(703) & cp_elements(713);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(711), clk => clk, reset => reset); --
    end block;
    rr_13231_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(711), ack => OR_u32_u32_3109_inst_req_0); -- 
    -- CP-element group 712 transition  output  bypass 
    -- predecessors 699 
    -- successors 715 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_3093_to_assign_stmt_3119/OR_u32_u32_3109_Update/cr
      -- 	branch_block_stmt_2042/assign_stmt_3093_to_assign_stmt_3119/OR_u32_u32_3109_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_3093_to_assign_stmt_3119/OR_u32_u32_3109_Update/$entry
      -- 
    cp_elements(712) <= cp_elements(699);
    cr_13236_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(712), ack => OR_u32_u32_3109_inst_req_1); -- 
    -- CP-element group 713 transition  bypass 
    -- predecessors 699 
    -- successors 711 
    -- members (4) 
      -- 	branch_block_stmt_2042/assign_stmt_3093_to_assign_stmt_3119/R_iNsTr_75_3108_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3093_to_assign_stmt_3119/R_iNsTr_75_3108_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_3093_to_assign_stmt_3119/R_iNsTr_75_3108_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3093_to_assign_stmt_3119/R_iNsTr_75_3108_sample_start_
      -- 
    cp_elements(713) <= cp_elements(699);
    -- CP-element group 714 transition  input  bypass 
    -- predecessors 711 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_3093_to_assign_stmt_3119/OR_u32_u32_3109_Sample/ra
      -- 	branch_block_stmt_2042/assign_stmt_3093_to_assign_stmt_3119/OR_u32_u32_3109_Sample/$exit
      -- 	branch_block_stmt_2042/assign_stmt_3093_to_assign_stmt_3119/OR_u32_u32_3109_sample_completed_
      -- 
    ra_13232_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => OR_u32_u32_3109_inst_ack_0, ack => cp_elements(714)); -- 
    -- CP-element group 715 transition  input  bypass 
    -- predecessors 712 
    -- successors 716 
    -- members (7) 
      -- 	branch_block_stmt_2042/assign_stmt_3093_to_assign_stmt_3119/OR_u32_u32_3109_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3093_to_assign_stmt_3119/R_iNsTr_132_3112_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3093_to_assign_stmt_3119/OR_u32_u32_3109_Update/$exit
      -- 	branch_block_stmt_2042/assign_stmt_3093_to_assign_stmt_3119/R_iNsTr_132_3112_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3093_to_assign_stmt_3119/R_iNsTr_132_3112_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_3093_to_assign_stmt_3119/R_iNsTr_132_3112_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_3093_to_assign_stmt_3119/OR_u32_u32_3109_Update/ca
      -- 
    ca_13237_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => OR_u32_u32_3109_inst_ack_1, ack => cp_elements(715)); -- 
    -- CP-element group 716 join  transition  output  bypass 
    -- predecessors 710 715 
    -- successors 718 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_3093_to_assign_stmt_3119/OR_u32_u32_3114_Sample/rr
      -- 	branch_block_stmt_2042/assign_stmt_3093_to_assign_stmt_3119/OR_u32_u32_3114_Sample/$entry
      -- 	branch_block_stmt_2042/assign_stmt_3093_to_assign_stmt_3119/OR_u32_u32_3114_sample_start_
      -- 
    cp_element_group_716: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 20) := "cp_element_group_716"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(710) & cp_elements(715);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(716), clk => clk, reset => reset); --
    end block;
    rr_13253_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(716), ack => OR_u32_u32_3114_inst_req_0); -- 
    -- CP-element group 717 transition  output  bypass 
    -- predecessors 699 
    -- successors 719 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_3093_to_assign_stmt_3119/OR_u32_u32_3114_Update/cr
      -- 	branch_block_stmt_2042/assign_stmt_3093_to_assign_stmt_3119/OR_u32_u32_3114_Update/$entry
      -- 	branch_block_stmt_2042/assign_stmt_3093_to_assign_stmt_3119/OR_u32_u32_3114_update_start_
      -- 
    cp_elements(717) <= cp_elements(699);
    cr_13258_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(717), ack => OR_u32_u32_3114_inst_req_1); -- 
    -- CP-element group 718 transition  input  bypass 
    -- predecessors 716 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_3093_to_assign_stmt_3119/OR_u32_u32_3114_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3093_to_assign_stmt_3119/OR_u32_u32_3114_Sample/ra
      -- 	branch_block_stmt_2042/assign_stmt_3093_to_assign_stmt_3119/OR_u32_u32_3114_Sample/$exit
      -- 
    ra_13254_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => OR_u32_u32_3114_inst_ack_0, ack => cp_elements(718)); -- 
    -- CP-element group 719 transition  input  output  bypass 
    -- predecessors 717 
    -- successors 721 
    -- members (10) 
      -- 	branch_block_stmt_2042/assign_stmt_3093_to_assign_stmt_3119/R_iNsTr_133_3117_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_3093_to_assign_stmt_3119/OR_u32_u32_3114_Update/ca
      -- 	branch_block_stmt_2042/assign_stmt_3093_to_assign_stmt_3119/OR_u32_u32_3114_Update/$exit
      -- 	branch_block_stmt_2042/assign_stmt_3093_to_assign_stmt_3119/R_iNsTr_133_3117_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3093_to_assign_stmt_3119/OR_u32_u32_3114_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3093_to_assign_stmt_3119/type_cast_3118_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_3093_to_assign_stmt_3119/R_iNsTr_133_3117_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3093_to_assign_stmt_3119/R_iNsTr_133_3117_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_3093_to_assign_stmt_3119/type_cast_3118_Sample/$entry
      -- 	branch_block_stmt_2042/assign_stmt_3093_to_assign_stmt_3119/type_cast_3118_Sample/rr
      -- 
    ca_13259_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => OR_u32_u32_3114_inst_ack_1, ack => cp_elements(719)); -- 
    rr_13271_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(719), ack => type_cast_3118_inst_req_0); -- 
    -- CP-element group 720 transition  output  bypass 
    -- predecessors 699 
    -- successors 722 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_3093_to_assign_stmt_3119/type_cast_3118_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_3093_to_assign_stmt_3119/type_cast_3118_Update/$entry
      -- 	branch_block_stmt_2042/assign_stmt_3093_to_assign_stmt_3119/type_cast_3118_Update/cr
      -- 
    cp_elements(720) <= cp_elements(699);
    cr_13276_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(720), ack => type_cast_3118_inst_req_1); -- 
    -- CP-element group 721 transition  input  bypass 
    -- predecessors 719 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_3093_to_assign_stmt_3119/type_cast_3118_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3093_to_assign_stmt_3119/type_cast_3118_Sample/$exit
      -- 	branch_block_stmt_2042/assign_stmt_3093_to_assign_stmt_3119/type_cast_3118_Sample/ra
      -- 
    ra_13272_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3118_inst_ack_0, ack => cp_elements(721)); -- 
    -- CP-element group 722 fork  transition  place  input  bypass 
    -- predecessors 720 
    -- successors 1974 1976 
    -- members (11) 
      -- 	branch_block_stmt_2042/assign_stmt_3093_to_assign_stmt_3119/type_cast_3118_update_completed_
      -- 	branch_block_stmt_2042/xx_xcritedgex_xix_xi28_omega_calcx_xexit
      -- 	branch_block_stmt_2042/assign_stmt_3093_to_assign_stmt_3119__exit__
      -- 	branch_block_stmt_2042/assign_stmt_3093_to_assign_stmt_3119/$exit
      -- 	branch_block_stmt_2042/assign_stmt_3093_to_assign_stmt_3119/type_cast_3118_Update/$exit
      -- 	branch_block_stmt_2042/assign_stmt_3093_to_assign_stmt_3119/type_cast_3118_Update/ca
      -- 	branch_block_stmt_2042/xx_xcritedgex_xix_xi28_omega_calcx_xexit_PhiReq/$entry
      -- 	branch_block_stmt_2042/xx_xcritedgex_xix_xi28_omega_calcx_xexit_PhiReq/phi_stmt_3122/$entry
      -- 	branch_block_stmt_2042/xx_xcritedgex_xix_xi28_omega_calcx_xexit_PhiReq/phi_stmt_3122/phi_stmt_3122_sources/$entry
      -- 	branch_block_stmt_2042/xx_xcritedgex_xix_xi28_omega_calcx_xexit_PhiReq/phi_stmt_3122/phi_stmt_3122_sources/type_cast_3125/$entry
      -- 	branch_block_stmt_2042/xx_xcritedgex_xix_xi28_omega_calcx_xexit_PhiReq/phi_stmt_3122/phi_stmt_3122_sources/type_cast_3125/SplitProtocol/$entry
      -- 
    ca_13277_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3118_inst_ack_1, ack => cp_elements(722)); -- 
    -- CP-element group 723 fork  transition  bypass 
    -- predecessors 1981 
    -- successors 724 725 728 729 732 733 736 740 743 744 
    -- members (1) 
      -- 	branch_block_stmt_2042/assign_stmt_3135_to_assign_stmt_3162/$entry
      -- 
    cp_elements(723) <= cp_elements(1981);
    -- CP-element group 724 transition  output  bypass 
    -- predecessors 723 
    -- successors 727 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_3135_to_assign_stmt_3162/SLT_f32_u1_3134_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_3135_to_assign_stmt_3162/SLT_f32_u1_3134_Update/$entry
      -- 	branch_block_stmt_2042/assign_stmt_3135_to_assign_stmt_3162/SLT_f32_u1_3134_Update/cr
      -- 
    cp_elements(724) <= cp_elements(723);
    cr_13297_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(724), ack => SLT_f32_u1_3134_inst_req_1); -- 
    -- CP-element group 725 transition  output  bypass 
    -- predecessors 723 
    -- successors 726 
    -- members (7) 
      -- 	branch_block_stmt_2042/assign_stmt_3135_to_assign_stmt_3162/SLT_f32_u1_3134_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_3135_to_assign_stmt_3162/R_iNsTr_42_3131_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_3135_to_assign_stmt_3162/R_iNsTr_42_3131_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3135_to_assign_stmt_3162/R_iNsTr_42_3131_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_3135_to_assign_stmt_3162/R_iNsTr_42_3131_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3135_to_assign_stmt_3162/SLT_f32_u1_3134_Sample/$entry
      -- 	branch_block_stmt_2042/assign_stmt_3135_to_assign_stmt_3162/SLT_f32_u1_3134_Sample/rr
      -- 
    cp_elements(725) <= cp_elements(723);
    rr_13292_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(725), ack => SLT_f32_u1_3134_inst_req_0); -- 
    -- CP-element group 726 transition  input  bypass 
    -- predecessors 725 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_3135_to_assign_stmt_3162/SLT_f32_u1_3134_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3135_to_assign_stmt_3162/SLT_f32_u1_3134_Sample/$exit
      -- 	branch_block_stmt_2042/assign_stmt_3135_to_assign_stmt_3162/SLT_f32_u1_3134_Sample/ra
      -- 
    ra_13293_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => SLT_f32_u1_3134_inst_ack_0, ack => cp_elements(726)); -- 
    -- CP-element group 727 transition  input  bypass 
    -- predecessors 724 
    -- successors 739 
    -- members (7) 
      -- 	branch_block_stmt_2042/assign_stmt_3135_to_assign_stmt_3162/SLT_f32_u1_3134_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3135_to_assign_stmt_3162/SLT_f32_u1_3134_Update/$exit
      -- 	branch_block_stmt_2042/assign_stmt_3135_to_assign_stmt_3162/SLT_f32_u1_3134_Update/ca
      -- 	branch_block_stmt_2042/assign_stmt_3135_to_assign_stmt_3162/R_iNsTr_60_3151_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_3135_to_assign_stmt_3162/R_iNsTr_60_3151_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3135_to_assign_stmt_3162/R_iNsTr_60_3151_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_3135_to_assign_stmt_3162/R_iNsTr_60_3151_update_completed_
      -- 
    ca_13298_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => SLT_f32_u1_3134_inst_ack_1, ack => cp_elements(727)); -- 
    -- CP-element group 728 transition  output  bypass 
    -- predecessors 723 
    -- successors 731 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_3135_to_assign_stmt_3162/MUL_f32_f32_3140_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_3135_to_assign_stmt_3162/MUL_f32_f32_3140_Update/$entry
      -- 	branch_block_stmt_2042/assign_stmt_3135_to_assign_stmt_3162/MUL_f32_f32_3140_Update/cr
      -- 
    cp_elements(728) <= cp_elements(723);
    cr_13315_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(728), ack => MUL_f32_f32_3140_inst_req_1); -- 
    -- CP-element group 729 transition  output  bypass 
    -- predecessors 723 
    -- successors 730 
    -- members (7) 
      -- 	branch_block_stmt_2042/assign_stmt_3135_to_assign_stmt_3162/MUL_f32_f32_3140_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_3135_to_assign_stmt_3162/R_iNsTr_42_3137_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_3135_to_assign_stmt_3162/R_iNsTr_42_3137_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3135_to_assign_stmt_3162/R_iNsTr_42_3137_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_3135_to_assign_stmt_3162/R_iNsTr_42_3137_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3135_to_assign_stmt_3162/MUL_f32_f32_3140_Sample/$entry
      -- 	branch_block_stmt_2042/assign_stmt_3135_to_assign_stmt_3162/MUL_f32_f32_3140_Sample/rr
      -- 
    cp_elements(729) <= cp_elements(723);
    rr_13310_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(729), ack => MUL_f32_f32_3140_inst_req_0); -- 
    -- CP-element group 730 transition  input  bypass 
    -- predecessors 729 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_3135_to_assign_stmt_3162/MUL_f32_f32_3140_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3135_to_assign_stmt_3162/MUL_f32_f32_3140_Sample/$exit
      -- 	branch_block_stmt_2042/assign_stmt_3135_to_assign_stmt_3162/MUL_f32_f32_3140_Sample/ra
      -- 
    ra_13311_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => MUL_f32_f32_3140_inst_ack_0, ack => cp_elements(730)); -- 
    -- CP-element group 731 transition  input  output  bypass 
    -- predecessors 728 
    -- successors 737 
    -- members (10) 
      -- 	branch_block_stmt_2042/assign_stmt_3135_to_assign_stmt_3162/MUL_f32_f32_3140_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3135_to_assign_stmt_3162/MUL_f32_f32_3140_Update/$exit
      -- 	branch_block_stmt_2042/assign_stmt_3135_to_assign_stmt_3162/MUL_f32_f32_3140_Update/ca
      -- 	branch_block_stmt_2042/assign_stmt_3135_to_assign_stmt_3162/type_cast_3148_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_3135_to_assign_stmt_3162/R_xx_xop_3147_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_3135_to_assign_stmt_3162/R_xx_xop_3147_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3135_to_assign_stmt_3162/R_xx_xop_3147_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_3135_to_assign_stmt_3162/R_xx_xop_3147_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3135_to_assign_stmt_3162/type_cast_3148_Sample/$entry
      -- 	branch_block_stmt_2042/assign_stmt_3135_to_assign_stmt_3162/type_cast_3148_Sample/rr
      -- 
    ca_13316_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => MUL_f32_f32_3140_inst_ack_1, ack => cp_elements(731)); -- 
    rr_13346_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(731), ack => type_cast_3148_inst_req_0); -- 
    -- CP-element group 732 transition  output  bypass 
    -- predecessors 723 
    -- successors 735 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_3135_to_assign_stmt_3162/type_cast_3144_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_3135_to_assign_stmt_3162/type_cast_3144_Update/$entry
      -- 	branch_block_stmt_2042/assign_stmt_3135_to_assign_stmt_3162/type_cast_3144_Update/cr
      -- 
    cp_elements(732) <= cp_elements(723);
    cr_13333_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(732), ack => type_cast_3144_inst_req_1); -- 
    -- CP-element group 733 transition  output  bypass 
    -- predecessors 723 
    -- successors 734 
    -- members (7) 
      -- 	branch_block_stmt_2042/assign_stmt_3135_to_assign_stmt_3162/type_cast_3144_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_3135_to_assign_stmt_3162/R_torque_refx_x0_3143_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_3135_to_assign_stmt_3162/R_torque_refx_x0_3143_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3135_to_assign_stmt_3162/R_torque_refx_x0_3143_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_3135_to_assign_stmt_3162/R_torque_refx_x0_3143_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3135_to_assign_stmt_3162/type_cast_3144_Sample/$entry
      -- 	branch_block_stmt_2042/assign_stmt_3135_to_assign_stmt_3162/type_cast_3144_Sample/rr
      -- 
    cp_elements(733) <= cp_elements(723);
    rr_13328_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(733), ack => type_cast_3144_inst_req_0); -- 
    -- CP-element group 734 transition  input  bypass 
    -- predecessors 733 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_3135_to_assign_stmt_3162/type_cast_3144_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3135_to_assign_stmt_3162/type_cast_3144_Sample/$exit
      -- 	branch_block_stmt_2042/assign_stmt_3135_to_assign_stmt_3162/type_cast_3144_Sample/ra
      -- 
    ra_13329_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3144_inst_ack_0, ack => cp_elements(734)); -- 
    -- CP-element group 735 transition  input  bypass 
    -- predecessors 732 
    -- successors 747 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_3135_to_assign_stmt_3162/type_cast_3144_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3135_to_assign_stmt_3162/type_cast_3144_Update/$exit
      -- 	branch_block_stmt_2042/assign_stmt_3135_to_assign_stmt_3162/type_cast_3144_Update/ca
      -- 
    ca_13334_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3144_inst_ack_1, ack => cp_elements(735)); -- 
    -- CP-element group 736 transition  output  bypass 
    -- predecessors 723 
    -- successors 738 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_3135_to_assign_stmt_3162/type_cast_3148_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_3135_to_assign_stmt_3162/type_cast_3148_Update/$entry
      -- 	branch_block_stmt_2042/assign_stmt_3135_to_assign_stmt_3162/type_cast_3148_Update/cr
      -- 
    cp_elements(736) <= cp_elements(723);
    cr_13351_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(736), ack => type_cast_3148_inst_req_1); -- 
    -- CP-element group 737 transition  input  bypass 
    -- predecessors 731 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_3135_to_assign_stmt_3162/type_cast_3148_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3135_to_assign_stmt_3162/type_cast_3148_Sample/$exit
      -- 	branch_block_stmt_2042/assign_stmt_3135_to_assign_stmt_3162/type_cast_3148_Sample/ra
      -- 
    ra_13347_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3148_inst_ack_0, ack => cp_elements(737)); -- 
    -- CP-element group 738 transition  input  bypass 
    -- predecessors 736 
    -- successors 739 
    -- members (7) 
      -- 	branch_block_stmt_2042/assign_stmt_3135_to_assign_stmt_3162/type_cast_3148_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3135_to_assign_stmt_3162/type_cast_3148_Update/$exit
      -- 	branch_block_stmt_2042/assign_stmt_3135_to_assign_stmt_3162/type_cast_3148_Update/ca
      -- 	branch_block_stmt_2042/assign_stmt_3135_to_assign_stmt_3162/R_iNsTr_61_3154_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_3135_to_assign_stmt_3162/R_iNsTr_61_3154_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3135_to_assign_stmt_3162/R_iNsTr_61_3154_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_3135_to_assign_stmt_3162/R_iNsTr_61_3154_update_completed_
      -- 
    ca_13352_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3148_inst_ack_1, ack => cp_elements(738)); -- 
    -- CP-element group 739 join  transition  output  bypass 
    -- predecessors 727 738 
    -- successors 741 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_3135_to_assign_stmt_3162/MUX_3155_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_3135_to_assign_stmt_3162/MUX_3155_start/$entry
      -- 	branch_block_stmt_2042/assign_stmt_3135_to_assign_stmt_3162/MUX_3155_start/req
      -- 
    cp_element_group_739: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 20) := "cp_element_group_739"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(727) & cp_elements(738);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(739), clk => clk, reset => reset); --
    end block;
    req_13368_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(739), ack => MUX_3155_inst_req_0); -- 
    -- CP-element group 740 transition  output  bypass 
    -- predecessors 723 
    -- successors 742 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_3135_to_assign_stmt_3162/MUX_3155_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_3135_to_assign_stmt_3162/MUX_3155_complete/$entry
      -- 	branch_block_stmt_2042/assign_stmt_3135_to_assign_stmt_3162/MUX_3155_complete/req
      -- 
    cp_elements(740) <= cp_elements(723);
    req_13373_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(740), ack => MUX_3155_inst_req_1); -- 
    -- CP-element group 741 transition  input  bypass 
    -- predecessors 739 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_3135_to_assign_stmt_3162/MUX_3155_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3135_to_assign_stmt_3162/MUX_3155_start/$exit
      -- 	branch_block_stmt_2042/assign_stmt_3135_to_assign_stmt_3162/MUX_3155_start/ack
      -- 
    ack_13369_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => MUX_3155_inst_ack_0, ack => cp_elements(741)); -- 
    -- CP-element group 742 transition  input  bypass 
    -- predecessors 740 
    -- successors 747 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_3135_to_assign_stmt_3162/MUX_3155_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3135_to_assign_stmt_3162/MUX_3155_complete/$exit
      -- 	branch_block_stmt_2042/assign_stmt_3135_to_assign_stmt_3162/MUX_3155_complete/ack
      -- 
    ack_13374_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => MUX_3155_inst_ack_1, ack => cp_elements(742)); -- 
    -- CP-element group 743 transition  output  bypass 
    -- predecessors 723 
    -- successors 746 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_3135_to_assign_stmt_3162/EQ_f32_u1_3161_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_3135_to_assign_stmt_3162/EQ_f32_u1_3161_Update/$entry
      -- 	branch_block_stmt_2042/assign_stmt_3135_to_assign_stmt_3162/EQ_f32_u1_3161_Update/cr
      -- 
    cp_elements(743) <= cp_elements(723);
    cr_13391_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(743), ack => EQ_f32_u1_3161_inst_req_1); -- 
    -- CP-element group 744 transition  output  bypass 
    -- predecessors 723 
    -- successors 745 
    -- members (7) 
      -- 	branch_block_stmt_2042/assign_stmt_3135_to_assign_stmt_3162/EQ_f32_u1_3161_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_3135_to_assign_stmt_3162/R_torque_refx_x0_3158_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_3135_to_assign_stmt_3162/R_torque_refx_x0_3158_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3135_to_assign_stmt_3162/R_torque_refx_x0_3158_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_3135_to_assign_stmt_3162/R_torque_refx_x0_3158_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3135_to_assign_stmt_3162/EQ_f32_u1_3161_Sample/$entry
      -- 	branch_block_stmt_2042/assign_stmt_3135_to_assign_stmt_3162/EQ_f32_u1_3161_Sample/rr
      -- 
    cp_elements(744) <= cp_elements(723);
    rr_13386_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(744), ack => EQ_f32_u1_3161_inst_req_0); -- 
    -- CP-element group 745 transition  input  bypass 
    -- predecessors 744 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_3135_to_assign_stmt_3162/EQ_f32_u1_3161_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3135_to_assign_stmt_3162/EQ_f32_u1_3161_Sample/$exit
      -- 	branch_block_stmt_2042/assign_stmt_3135_to_assign_stmt_3162/EQ_f32_u1_3161_Sample/ra
      -- 
    ra_13387_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_f32_u1_3161_inst_ack_0, ack => cp_elements(745)); -- 
    -- CP-element group 746 transition  input  bypass 
    -- predecessors 743 
    -- successors 747 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_3135_to_assign_stmt_3162/EQ_f32_u1_3161_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3135_to_assign_stmt_3162/EQ_f32_u1_3161_Update/$exit
      -- 	branch_block_stmt_2042/assign_stmt_3135_to_assign_stmt_3162/EQ_f32_u1_3161_Update/ca
      -- 
    ca_13392_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_f32_u1_3161_inst_ack_1, ack => cp_elements(746)); -- 
    -- CP-element group 747 join  transition  bypass 
    -- predecessors 735 742 746 
    -- successors 43 
    -- members (1) 
      -- 	branch_block_stmt_2042/assign_stmt_3135_to_assign_stmt_3162/$exit
      -- 
    cp_element_group_747: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 20) := "cp_element_group_747"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= cp_elements(735) & cp_elements(742) & cp_elements(746);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(747), clk => clk, reset => reset); --
    end block;
    -- CP-element group 748 transition  place  dead  bypass 
    -- predecessors 43 
    -- successors 44 
    -- members (8) 
      -- 	branch_block_stmt_2042/merge_stmt_3169__entry__
      -- 	branch_block_stmt_2042/if_stmt_3163__exit__
      -- 	branch_block_stmt_2042/if_stmt_3163_dead_link/$entry
      -- 	branch_block_stmt_2042/if_stmt_3163_dead_link/$exit
      -- 	branch_block_stmt_2042/if_stmt_3163_dead_link/dead_transition
      -- 	branch_block_stmt_2042/merge_stmt_3169_dead_link/$entry
      -- 	branch_block_stmt_2042/merge_stmt_3169_dead_link/$exit
      -- 	branch_block_stmt_2042/merge_stmt_3169_dead_link/dead_transition
      -- 
    cp_elements(748) <= false;
    -- CP-element group 749 transition  output  bypass 
    -- predecessors 43 
    -- successors 750 
    -- members (3) 
      -- 	branch_block_stmt_2042/if_stmt_3163_eval_test/$entry
      -- 	branch_block_stmt_2042/if_stmt_3163_eval_test/$exit
      -- 	branch_block_stmt_2042/if_stmt_3163_eval_test/branch_req
      -- 
    cp_elements(749) <= cp_elements(43);
    branch_req_13400_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(749), ack => if_stmt_3163_branch_req_0); -- 
    -- CP-element group 750 branch  place  bypass 
    -- predecessors 749 
    -- successors 751 753 
    -- members (1) 
      -- 	branch_block_stmt_2042/R_iNsTr_62_3164_place
      -- 
    cp_elements(750) <= cp_elements(749);
    -- CP-element group 751 transition  bypass 
    -- predecessors 750 
    -- successors 752 
    -- members (1) 
      -- 	branch_block_stmt_2042/if_stmt_3163_if_link/$entry
      -- 
    cp_elements(751) <= cp_elements(750);
    -- CP-element group 752 fork  transition  place  input  bypass 
    -- predecessors 751 
    -- successors 2291 2292 
    -- members (8) 
      -- 	branch_block_stmt_2042/omega_calcx_xexit_iq_err_calcx_xexit
      -- 	branch_block_stmt_2042/if_stmt_3163_if_link/$exit
      -- 	branch_block_stmt_2042/if_stmt_3163_if_link/if_choice_transition
      -- 	branch_block_stmt_2042/omega_calcx_xexit_iq_err_calcx_xexit_PhiReq/$entry
      -- 	branch_block_stmt_2042/omega_calcx_xexit_iq_err_calcx_xexit_PhiReq/phi_stmt_3568/$entry
      -- 	branch_block_stmt_2042/omega_calcx_xexit_iq_err_calcx_xexit_PhiReq/phi_stmt_3568/phi_stmt_3568_sources/$entry
      -- 	branch_block_stmt_2042/omega_calcx_xexit_iq_err_calcx_xexit_PhiReq/phi_stmt_3568/phi_stmt_3568_sources/type_cast_3571/$entry
      -- 	branch_block_stmt_2042/omega_calcx_xexit_iq_err_calcx_xexit_PhiReq/phi_stmt_3568/phi_stmt_3568_sources/type_cast_3571/SplitProtocol/$entry
      -- 
    if_choice_transition_13405_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_3163_branch_ack_1, ack => cp_elements(752)); -- 
    -- CP-element group 753 transition  bypass 
    -- predecessors 750 
    -- successors 754 
    -- members (1) 
      -- 	branch_block_stmt_2042/if_stmt_3163_else_link/$entry
      -- 
    cp_elements(753) <= cp_elements(750);
    -- CP-element group 754 transition  place  input  bypass 
    -- predecessors 753 
    -- successors 44 
    -- members (9) 
      -- 	branch_block_stmt_2042/omega_calcx_xexit_bb_41
      -- 	branch_block_stmt_2042/if_stmt_3163_else_link/$exit
      -- 	branch_block_stmt_2042/if_stmt_3163_else_link/else_choice_transition
      -- 	branch_block_stmt_2042/merge_stmt_3169_PhiReqMerge
      -- 	branch_block_stmt_2042/omega_calcx_xexit_bb_41_PhiReq/$entry
      -- 	branch_block_stmt_2042/omega_calcx_xexit_bb_41_PhiReq/$exit
      -- 	branch_block_stmt_2042/merge_stmt_3169_PhiAck/$entry
      -- 	branch_block_stmt_2042/merge_stmt_3169_PhiAck/$exit
      -- 	branch_block_stmt_2042/merge_stmt_3169_PhiAck/dummy
      -- 
    else_choice_transition_13409_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_3163_branch_ack_0, ack => cp_elements(754)); -- 
    -- CP-element group 755 fork  transition  bypass 
    -- predecessors 44 
    -- successors 756 757 760 763 764 767 770 771 774 777 780 781 784 787 791 792 793 796 800 
    -- members (1) 
      -- 	branch_block_stmt_2042/assign_stmt_3175_to_assign_stmt_3245/$entry
      -- 
    cp_elements(755) <= cp_elements(44);
    -- CP-element group 756 transition  output  bypass 
    -- predecessors 755 
    -- successors 759 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_3175_to_assign_stmt_3245/LSHR_u32_u32_3174_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_3175_to_assign_stmt_3245/LSHR_u32_u32_3174_Update/$entry
      -- 	branch_block_stmt_2042/assign_stmt_3175_to_assign_stmt_3245/LSHR_u32_u32_3174_Update/cr
      -- 
    cp_elements(756) <= cp_elements(755);
    cr_13431_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(756), ack => LSHR_u32_u32_3174_inst_req_1); -- 
    -- CP-element group 757 transition  output  bypass 
    -- predecessors 755 
    -- successors 758 
    -- members (7) 
      -- 	branch_block_stmt_2042/assign_stmt_3175_to_assign_stmt_3245/LSHR_u32_u32_3174_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_3175_to_assign_stmt_3245/R_tmp10x_xix_xi_3171_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_3175_to_assign_stmt_3245/R_tmp10x_xix_xi_3171_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3175_to_assign_stmt_3245/R_tmp10x_xix_xi_3171_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_3175_to_assign_stmt_3245/R_tmp10x_xix_xi_3171_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3175_to_assign_stmt_3245/LSHR_u32_u32_3174_Sample/$entry
      -- 	branch_block_stmt_2042/assign_stmt_3175_to_assign_stmt_3245/LSHR_u32_u32_3174_Sample/rr
      -- 
    cp_elements(757) <= cp_elements(755);
    rr_13426_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(757), ack => LSHR_u32_u32_3174_inst_req_0); -- 
    -- CP-element group 758 transition  input  bypass 
    -- predecessors 757 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_3175_to_assign_stmt_3245/LSHR_u32_u32_3174_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3175_to_assign_stmt_3245/LSHR_u32_u32_3174_Sample/$exit
      -- 	branch_block_stmt_2042/assign_stmt_3175_to_assign_stmt_3245/LSHR_u32_u32_3174_Sample/ra
      -- 
    ra_13427_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => LSHR_u32_u32_3174_inst_ack_0, ack => cp_elements(758)); -- 
    -- CP-element group 759 transition  input  output  bypass 
    -- predecessors 756 
    -- successors 761 
    -- members (10) 
      -- 	branch_block_stmt_2042/assign_stmt_3175_to_assign_stmt_3245/LSHR_u32_u32_3174_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3175_to_assign_stmt_3245/LSHR_u32_u32_3174_Update/$exit
      -- 	branch_block_stmt_2042/assign_stmt_3175_to_assign_stmt_3245/LSHR_u32_u32_3174_Update/ca
      -- 	branch_block_stmt_2042/assign_stmt_3175_to_assign_stmt_3245/AND_u32_u32_3180_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_3175_to_assign_stmt_3245/R_iNsTr_88_3177_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_3175_to_assign_stmt_3245/R_iNsTr_88_3177_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3175_to_assign_stmt_3245/R_iNsTr_88_3177_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_3175_to_assign_stmt_3245/R_iNsTr_88_3177_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3175_to_assign_stmt_3245/AND_u32_u32_3180_Sample/$entry
      -- 	branch_block_stmt_2042/assign_stmt_3175_to_assign_stmt_3245/AND_u32_u32_3180_Sample/rr
      -- 
    ca_13432_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => LSHR_u32_u32_3174_inst_ack_1, ack => cp_elements(759)); -- 
    rr_13444_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(759), ack => AND_u32_u32_3180_inst_req_0); -- 
    -- CP-element group 760 transition  output  bypass 
    -- predecessors 755 
    -- successors 762 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_3175_to_assign_stmt_3245/AND_u32_u32_3180_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_3175_to_assign_stmt_3245/AND_u32_u32_3180_Update/$entry
      -- 	branch_block_stmt_2042/assign_stmt_3175_to_assign_stmt_3245/AND_u32_u32_3180_Update/cr
      -- 
    cp_elements(760) <= cp_elements(755);
    cr_13449_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(760), ack => AND_u32_u32_3180_inst_req_1); -- 
    -- CP-element group 761 transition  input  bypass 
    -- predecessors 759 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_3175_to_assign_stmt_3245/AND_u32_u32_3180_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3175_to_assign_stmt_3245/AND_u32_u32_3180_Sample/$exit
      -- 	branch_block_stmt_2042/assign_stmt_3175_to_assign_stmt_3245/AND_u32_u32_3180_Sample/ra
      -- 
    ra_13445_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => AND_u32_u32_3180_inst_ack_0, ack => cp_elements(761)); -- 
    -- CP-element group 762 transition  input  bypass 
    -- predecessors 760 
    -- successors 799 
    -- members (7) 
      -- 	branch_block_stmt_2042/assign_stmt_3175_to_assign_stmt_3245/AND_u32_u32_3180_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3175_to_assign_stmt_3245/AND_u32_u32_3180_Update/$exit
      -- 	branch_block_stmt_2042/assign_stmt_3175_to_assign_stmt_3245/AND_u32_u32_3180_Update/ca
      -- 	branch_block_stmt_2042/assign_stmt_3175_to_assign_stmt_3245/R_iNsTr_89_3242_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3175_to_assign_stmt_3245/R_iNsTr_89_3242_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_3175_to_assign_stmt_3245/R_iNsTr_89_3242_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_3175_to_assign_stmt_3245/R_iNsTr_89_3242_update_completed_
      -- 
    ca_13450_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => AND_u32_u32_3180_inst_ack_1, ack => cp_elements(762)); -- 
    -- CP-element group 763 transition  output  bypass 
    -- predecessors 755 
    -- successors 766 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_3175_to_assign_stmt_3245/LSHR_u32_u32_3186_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_3175_to_assign_stmt_3245/LSHR_u32_u32_3186_Update/$entry
      -- 	branch_block_stmt_2042/assign_stmt_3175_to_assign_stmt_3245/LSHR_u32_u32_3186_Update/cr
      -- 
    cp_elements(763) <= cp_elements(755);
    cr_13467_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(763), ack => LSHR_u32_u32_3186_inst_req_1); -- 
    -- CP-element group 764 transition  output  bypass 
    -- predecessors 755 
    -- successors 765 
    -- members (7) 
      -- 	branch_block_stmt_2042/assign_stmt_3175_to_assign_stmt_3245/LSHR_u32_u32_3186_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_3175_to_assign_stmt_3245/R_tmp6x_xix_xi_3183_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_3175_to_assign_stmt_3245/R_tmp6x_xix_xi_3183_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3175_to_assign_stmt_3245/R_tmp6x_xix_xi_3183_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_3175_to_assign_stmt_3245/R_tmp6x_xix_xi_3183_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3175_to_assign_stmt_3245/LSHR_u32_u32_3186_Sample/$entry
      -- 	branch_block_stmt_2042/assign_stmt_3175_to_assign_stmt_3245/LSHR_u32_u32_3186_Sample/rr
      -- 
    cp_elements(764) <= cp_elements(755);
    rr_13462_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(764), ack => LSHR_u32_u32_3186_inst_req_0); -- 
    -- CP-element group 765 transition  input  bypass 
    -- predecessors 764 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_3175_to_assign_stmt_3245/LSHR_u32_u32_3186_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3175_to_assign_stmt_3245/LSHR_u32_u32_3186_Sample/$exit
      -- 	branch_block_stmt_2042/assign_stmt_3175_to_assign_stmt_3245/LSHR_u32_u32_3186_Sample/ra
      -- 
    ra_13463_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => LSHR_u32_u32_3186_inst_ack_0, ack => cp_elements(765)); -- 
    -- CP-element group 766 transition  input  output  bypass 
    -- predecessors 763 
    -- successors 768 
    -- members (10) 
      -- 	branch_block_stmt_2042/assign_stmt_3175_to_assign_stmt_3245/LSHR_u32_u32_3186_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3175_to_assign_stmt_3245/LSHR_u32_u32_3186_Update/$exit
      -- 	branch_block_stmt_2042/assign_stmt_3175_to_assign_stmt_3245/LSHR_u32_u32_3186_Update/ca
      -- 	branch_block_stmt_2042/assign_stmt_3175_to_assign_stmt_3245/AND_u32_u32_3192_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_3175_to_assign_stmt_3245/R_iNsTr_90_3189_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_3175_to_assign_stmt_3245/R_iNsTr_90_3189_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3175_to_assign_stmt_3245/R_iNsTr_90_3189_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_3175_to_assign_stmt_3245/R_iNsTr_90_3189_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3175_to_assign_stmt_3245/AND_u32_u32_3192_Sample/$entry
      -- 	branch_block_stmt_2042/assign_stmt_3175_to_assign_stmt_3245/AND_u32_u32_3192_Sample/rr
      -- 
    ca_13468_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => LSHR_u32_u32_3186_inst_ack_1, ack => cp_elements(766)); -- 
    rr_13480_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(766), ack => AND_u32_u32_3192_inst_req_0); -- 
    -- CP-element group 767 transition  output  bypass 
    -- predecessors 755 
    -- successors 769 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_3175_to_assign_stmt_3245/AND_u32_u32_3192_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_3175_to_assign_stmt_3245/AND_u32_u32_3192_Update/$entry
      -- 	branch_block_stmt_2042/assign_stmt_3175_to_assign_stmt_3245/AND_u32_u32_3192_Update/cr
      -- 
    cp_elements(767) <= cp_elements(755);
    cr_13485_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(767), ack => AND_u32_u32_3192_inst_req_1); -- 
    -- CP-element group 768 transition  input  bypass 
    -- predecessors 766 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_3175_to_assign_stmt_3245/AND_u32_u32_3192_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3175_to_assign_stmt_3245/AND_u32_u32_3192_Sample/$exit
      -- 	branch_block_stmt_2042/assign_stmt_3175_to_assign_stmt_3245/AND_u32_u32_3192_Sample/ra
      -- 
    ra_13481_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => AND_u32_u32_3192_inst_ack_0, ack => cp_elements(768)); -- 
    -- CP-element group 769 transition  input  bypass 
    -- predecessors 767 
    -- successors 799 
    -- members (7) 
      -- 	branch_block_stmt_2042/assign_stmt_3175_to_assign_stmt_3245/AND_u32_u32_3192_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3175_to_assign_stmt_3245/AND_u32_u32_3192_Update/$exit
      -- 	branch_block_stmt_2042/assign_stmt_3175_to_assign_stmt_3245/AND_u32_u32_3192_Update/ca
      -- 	branch_block_stmt_2042/assign_stmt_3175_to_assign_stmt_3245/R_iNsTr_91_3243_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_3175_to_assign_stmt_3245/R_iNsTr_91_3243_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3175_to_assign_stmt_3245/R_iNsTr_91_3243_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_3175_to_assign_stmt_3245/R_iNsTr_91_3243_update_completed_
      -- 
    ca_13486_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => AND_u32_u32_3192_inst_ack_1, ack => cp_elements(769)); -- 
    -- CP-element group 770 transition  output  bypass 
    -- predecessors 755 
    -- successors 773 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_3175_to_assign_stmt_3245/SHL_u32_u32_3198_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_3175_to_assign_stmt_3245/SHL_u32_u32_3198_Update/$entry
      -- 	branch_block_stmt_2042/assign_stmt_3175_to_assign_stmt_3245/SHL_u32_u32_3198_Update/cr
      -- 
    cp_elements(770) <= cp_elements(755);
    cr_13503_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(770), ack => SHL_u32_u32_3198_inst_req_1); -- 
    -- CP-element group 771 transition  output  bypass 
    -- predecessors 755 
    -- successors 772 
    -- members (7) 
      -- 	branch_block_stmt_2042/assign_stmt_3175_to_assign_stmt_3245/SHL_u32_u32_3198_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_3175_to_assign_stmt_3245/R_tmp10x_xix_xi_3195_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_3175_to_assign_stmt_3245/R_tmp10x_xix_xi_3195_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3175_to_assign_stmt_3245/R_tmp10x_xix_xi_3195_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_3175_to_assign_stmt_3245/R_tmp10x_xix_xi_3195_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3175_to_assign_stmt_3245/SHL_u32_u32_3198_Sample/$entry
      -- 	branch_block_stmt_2042/assign_stmt_3175_to_assign_stmt_3245/SHL_u32_u32_3198_Sample/rr
      -- 
    cp_elements(771) <= cp_elements(755);
    rr_13498_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(771), ack => SHL_u32_u32_3198_inst_req_0); -- 
    -- CP-element group 772 transition  input  bypass 
    -- predecessors 771 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_3175_to_assign_stmt_3245/SHL_u32_u32_3198_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3175_to_assign_stmt_3245/SHL_u32_u32_3198_Sample/$exit
      -- 	branch_block_stmt_2042/assign_stmt_3175_to_assign_stmt_3245/SHL_u32_u32_3198_Sample/ra
      -- 
    ra_13499_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => SHL_u32_u32_3198_inst_ack_0, ack => cp_elements(772)); -- 
    -- CP-element group 773 transition  input  output  bypass 
    -- predecessors 770 
    -- successors 775 
    -- members (10) 
      -- 	branch_block_stmt_2042/assign_stmt_3175_to_assign_stmt_3245/SHL_u32_u32_3198_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3175_to_assign_stmt_3245/SHL_u32_u32_3198_Update/$exit
      -- 	branch_block_stmt_2042/assign_stmt_3175_to_assign_stmt_3245/SHL_u32_u32_3198_Update/ca
      -- 	branch_block_stmt_2042/assign_stmt_3175_to_assign_stmt_3245/AND_u32_u32_3204_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_3175_to_assign_stmt_3245/R_iNsTr_92_3201_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_3175_to_assign_stmt_3245/R_iNsTr_92_3201_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3175_to_assign_stmt_3245/R_iNsTr_92_3201_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_3175_to_assign_stmt_3245/R_iNsTr_92_3201_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3175_to_assign_stmt_3245/AND_u32_u32_3204_Sample/$entry
      -- 	branch_block_stmt_2042/assign_stmt_3175_to_assign_stmt_3245/AND_u32_u32_3204_Sample/rr
      -- 
    ca_13504_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => SHL_u32_u32_3198_inst_ack_1, ack => cp_elements(773)); -- 
    rr_13516_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(773), ack => AND_u32_u32_3204_inst_req_0); -- 
    -- CP-element group 774 transition  output  bypass 
    -- predecessors 755 
    -- successors 776 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_3175_to_assign_stmt_3245/AND_u32_u32_3204_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_3175_to_assign_stmt_3245/AND_u32_u32_3204_Update/$entry
      -- 	branch_block_stmt_2042/assign_stmt_3175_to_assign_stmt_3245/AND_u32_u32_3204_Update/cr
      -- 
    cp_elements(774) <= cp_elements(755);
    cr_13521_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(774), ack => AND_u32_u32_3204_inst_req_1); -- 
    -- CP-element group 775 transition  input  bypass 
    -- predecessors 773 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_3175_to_assign_stmt_3245/AND_u32_u32_3204_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3175_to_assign_stmt_3245/AND_u32_u32_3204_Sample/$exit
      -- 	branch_block_stmt_2042/assign_stmt_3175_to_assign_stmt_3245/AND_u32_u32_3204_Sample/ra
      -- 
    ra_13517_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => AND_u32_u32_3204_inst_ack_0, ack => cp_elements(775)); -- 
    -- CP-element group 776 transition  input  output  bypass 
    -- predecessors 774 
    -- successors 778 
    -- members (10) 
      -- 	branch_block_stmt_2042/assign_stmt_3175_to_assign_stmt_3245/AND_u32_u32_3204_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3175_to_assign_stmt_3245/AND_u32_u32_3204_Update/$exit
      -- 	branch_block_stmt_2042/assign_stmt_3175_to_assign_stmt_3245/AND_u32_u32_3204_Update/ca
      -- 	branch_block_stmt_2042/assign_stmt_3175_to_assign_stmt_3245/OR_u32_u32_3210_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_3175_to_assign_stmt_3245/R_iNsTr_93_3207_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_3175_to_assign_stmt_3245/R_iNsTr_93_3207_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3175_to_assign_stmt_3245/R_iNsTr_93_3207_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_3175_to_assign_stmt_3245/R_iNsTr_93_3207_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3175_to_assign_stmt_3245/OR_u32_u32_3210_Sample/$entry
      -- 	branch_block_stmt_2042/assign_stmt_3175_to_assign_stmt_3245/OR_u32_u32_3210_Sample/rr
      -- 
    ca_13522_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => AND_u32_u32_3204_inst_ack_1, ack => cp_elements(776)); -- 
    rr_13534_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(776), ack => OR_u32_u32_3210_inst_req_0); -- 
    -- CP-element group 777 transition  output  bypass 
    -- predecessors 755 
    -- successors 779 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_3175_to_assign_stmt_3245/OR_u32_u32_3210_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_3175_to_assign_stmt_3245/OR_u32_u32_3210_Update/$entry
      -- 	branch_block_stmt_2042/assign_stmt_3175_to_assign_stmt_3245/OR_u32_u32_3210_Update/cr
      -- 
    cp_elements(777) <= cp_elements(755);
    cr_13539_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(777), ack => OR_u32_u32_3210_inst_req_1); -- 
    -- CP-element group 778 transition  input  bypass 
    -- predecessors 776 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_3175_to_assign_stmt_3245/OR_u32_u32_3210_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3175_to_assign_stmt_3245/OR_u32_u32_3210_Sample/$exit
      -- 	branch_block_stmt_2042/assign_stmt_3175_to_assign_stmt_3245/OR_u32_u32_3210_Sample/ra
      -- 
    ra_13535_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => OR_u32_u32_3210_inst_ack_0, ack => cp_elements(778)); -- 
    -- CP-element group 779 transition  input  bypass 
    -- predecessors 777 
    -- successors 803 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_3175_to_assign_stmt_3245/OR_u32_u32_3210_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3175_to_assign_stmt_3245/OR_u32_u32_3210_Update/$exit
      -- 	branch_block_stmt_2042/assign_stmt_3175_to_assign_stmt_3245/OR_u32_u32_3210_Update/ca
      -- 
    ca_13540_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => OR_u32_u32_3210_inst_ack_1, ack => cp_elements(779)); -- 
    -- CP-element group 780 transition  output  bypass 
    -- predecessors 755 
    -- successors 783 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_3175_to_assign_stmt_3245/LSHR_u32_u32_3216_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_3175_to_assign_stmt_3245/LSHR_u32_u32_3216_Update/$entry
      -- 	branch_block_stmt_2042/assign_stmt_3175_to_assign_stmt_3245/LSHR_u32_u32_3216_Update/cr
      -- 
    cp_elements(780) <= cp_elements(755);
    cr_13557_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(780), ack => LSHR_u32_u32_3216_inst_req_1); -- 
    -- CP-element group 781 transition  output  bypass 
    -- predecessors 755 
    -- successors 782 
    -- members (7) 
      -- 	branch_block_stmt_2042/assign_stmt_3175_to_assign_stmt_3245/LSHR_u32_u32_3216_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_3175_to_assign_stmt_3245/R_tmp6x_xix_xi_3213_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_3175_to_assign_stmt_3245/R_tmp6x_xix_xi_3213_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3175_to_assign_stmt_3245/R_tmp6x_xix_xi_3213_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_3175_to_assign_stmt_3245/R_tmp6x_xix_xi_3213_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3175_to_assign_stmt_3245/LSHR_u32_u32_3216_Sample/$entry
      -- 	branch_block_stmt_2042/assign_stmt_3175_to_assign_stmt_3245/LSHR_u32_u32_3216_Sample/rr
      -- 
    cp_elements(781) <= cp_elements(755);
    rr_13552_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(781), ack => LSHR_u32_u32_3216_inst_req_0); -- 
    -- CP-element group 782 transition  input  bypass 
    -- predecessors 781 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_3175_to_assign_stmt_3245/LSHR_u32_u32_3216_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3175_to_assign_stmt_3245/LSHR_u32_u32_3216_Sample/$exit
      -- 	branch_block_stmt_2042/assign_stmt_3175_to_assign_stmt_3245/LSHR_u32_u32_3216_Sample/ra
      -- 
    ra_13553_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => LSHR_u32_u32_3216_inst_ack_0, ack => cp_elements(782)); -- 
    -- CP-element group 783 transition  input  output  bypass 
    -- predecessors 780 
    -- successors 785 
    -- members (10) 
      -- 	branch_block_stmt_2042/assign_stmt_3175_to_assign_stmt_3245/LSHR_u32_u32_3216_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3175_to_assign_stmt_3245/LSHR_u32_u32_3216_Update/$exit
      -- 	branch_block_stmt_2042/assign_stmt_3175_to_assign_stmt_3245/LSHR_u32_u32_3216_Update/ca
      -- 	branch_block_stmt_2042/assign_stmt_3175_to_assign_stmt_3245/AND_u32_u32_3222_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_3175_to_assign_stmt_3245/R_iNsTr_95_3219_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_3175_to_assign_stmt_3245/R_iNsTr_95_3219_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3175_to_assign_stmt_3245/R_iNsTr_95_3219_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_3175_to_assign_stmt_3245/R_iNsTr_95_3219_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3175_to_assign_stmt_3245/AND_u32_u32_3222_Sample/$entry
      -- 	branch_block_stmt_2042/assign_stmt_3175_to_assign_stmt_3245/AND_u32_u32_3222_Sample/rr
      -- 
    ca_13558_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => LSHR_u32_u32_3216_inst_ack_1, ack => cp_elements(783)); -- 
    rr_13570_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(783), ack => AND_u32_u32_3222_inst_req_0); -- 
    -- CP-element group 784 transition  output  bypass 
    -- predecessors 755 
    -- successors 786 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_3175_to_assign_stmt_3245/AND_u32_u32_3222_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_3175_to_assign_stmt_3245/AND_u32_u32_3222_Update/$entry
      -- 	branch_block_stmt_2042/assign_stmt_3175_to_assign_stmt_3245/AND_u32_u32_3222_Update/cr
      -- 
    cp_elements(784) <= cp_elements(755);
    cr_13575_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(784), ack => AND_u32_u32_3222_inst_req_1); -- 
    -- CP-element group 785 transition  input  bypass 
    -- predecessors 783 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_3175_to_assign_stmt_3245/AND_u32_u32_3222_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3175_to_assign_stmt_3245/AND_u32_u32_3222_Sample/$exit
      -- 	branch_block_stmt_2042/assign_stmt_3175_to_assign_stmt_3245/AND_u32_u32_3222_Sample/ra
      -- 
    ra_13571_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => AND_u32_u32_3222_inst_ack_0, ack => cp_elements(785)); -- 
    -- CP-element group 786 transition  input  output  bypass 
    -- predecessors 784 
    -- successors 788 
    -- members (10) 
      -- 	branch_block_stmt_2042/assign_stmt_3175_to_assign_stmt_3245/AND_u32_u32_3222_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3175_to_assign_stmt_3245/AND_u32_u32_3222_Update/$exit
      -- 	branch_block_stmt_2042/assign_stmt_3175_to_assign_stmt_3245/AND_u32_u32_3222_Update/ca
      -- 	branch_block_stmt_2042/assign_stmt_3175_to_assign_stmt_3245/OR_u32_u32_3228_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_3175_to_assign_stmt_3245/R_iNsTr_96_3225_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_3175_to_assign_stmt_3245/R_iNsTr_96_3225_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3175_to_assign_stmt_3245/R_iNsTr_96_3225_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_3175_to_assign_stmt_3245/R_iNsTr_96_3225_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3175_to_assign_stmt_3245/OR_u32_u32_3228_Sample/$entry
      -- 	branch_block_stmt_2042/assign_stmt_3175_to_assign_stmt_3245/OR_u32_u32_3228_Sample/rr
      -- 
    ca_13576_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => AND_u32_u32_3222_inst_ack_1, ack => cp_elements(786)); -- 
    rr_13588_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(786), ack => OR_u32_u32_3228_inst_req_0); -- 
    -- CP-element group 787 transition  output  bypass 
    -- predecessors 755 
    -- successors 789 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_3175_to_assign_stmt_3245/OR_u32_u32_3228_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_3175_to_assign_stmt_3245/OR_u32_u32_3228_Update/$entry
      -- 	branch_block_stmt_2042/assign_stmt_3175_to_assign_stmt_3245/OR_u32_u32_3228_Update/cr
      -- 
    cp_elements(787) <= cp_elements(755);
    cr_13593_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(787), ack => OR_u32_u32_3228_inst_req_1); -- 
    -- CP-element group 788 transition  input  bypass 
    -- predecessors 786 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_3175_to_assign_stmt_3245/OR_u32_u32_3228_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3175_to_assign_stmt_3245/OR_u32_u32_3228_Sample/$exit
      -- 	branch_block_stmt_2042/assign_stmt_3175_to_assign_stmt_3245/OR_u32_u32_3228_Sample/ra
      -- 
    ra_13589_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => OR_u32_u32_3228_inst_ack_0, ack => cp_elements(788)); -- 
    -- CP-element group 789 transition  input  bypass 
    -- predecessors 787 
    -- successors 803 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_3175_to_assign_stmt_3245/OR_u32_u32_3228_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3175_to_assign_stmt_3245/OR_u32_u32_3228_Update/$exit
      -- 	branch_block_stmt_2042/assign_stmt_3175_to_assign_stmt_3245/OR_u32_u32_3228_Update/ca
      -- 
    ca_13594_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => OR_u32_u32_3228_inst_ack_1, ack => cp_elements(789)); -- 
    -- CP-element group 790 join  transition  output  bypass 
    -- predecessors 792 793 
    -- successors 794 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_3175_to_assign_stmt_3245/XOR_u32_u32_3233_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_3175_to_assign_stmt_3245/XOR_u32_u32_3233_Sample/$entry
      -- 	branch_block_stmt_2042/assign_stmt_3175_to_assign_stmt_3245/XOR_u32_u32_3233_Sample/rr
      -- 
    cp_element_group_790: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 20) := "cp_element_group_790"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(792) & cp_elements(793);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(790), clk => clk, reset => reset); --
    end block;
    rr_13610_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(790), ack => XOR_u32_u32_3233_inst_req_0); -- 
    -- CP-element group 791 transition  output  bypass 
    -- predecessors 755 
    -- successors 795 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_3175_to_assign_stmt_3245/XOR_u32_u32_3233_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_3175_to_assign_stmt_3245/XOR_u32_u32_3233_Update/$entry
      -- 	branch_block_stmt_2042/assign_stmt_3175_to_assign_stmt_3245/XOR_u32_u32_3233_Update/cr
      -- 
    cp_elements(791) <= cp_elements(755);
    cr_13615_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(791), ack => XOR_u32_u32_3233_inst_req_1); -- 
    -- CP-element group 792 transition  bypass 
    -- predecessors 755 
    -- successors 790 
    -- members (4) 
      -- 	branch_block_stmt_2042/assign_stmt_3175_to_assign_stmt_3245/R_tmp6x_xix_xi_3231_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_3175_to_assign_stmt_3245/R_tmp6x_xix_xi_3231_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3175_to_assign_stmt_3245/R_tmp6x_xix_xi_3231_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_3175_to_assign_stmt_3245/R_tmp6x_xix_xi_3231_update_completed_
      -- 
    cp_elements(792) <= cp_elements(755);
    -- CP-element group 793 transition  bypass 
    -- predecessors 755 
    -- successors 790 
    -- members (4) 
      -- 	branch_block_stmt_2042/assign_stmt_3175_to_assign_stmt_3245/R_tmp10x_xix_xi_3232_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_3175_to_assign_stmt_3245/R_tmp10x_xix_xi_3232_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3175_to_assign_stmt_3245/R_tmp10x_xix_xi_3232_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_3175_to_assign_stmt_3245/R_tmp10x_xix_xi_3232_update_completed_
      -- 
    cp_elements(793) <= cp_elements(755);
    -- CP-element group 794 transition  input  bypass 
    -- predecessors 790 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_3175_to_assign_stmt_3245/XOR_u32_u32_3233_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3175_to_assign_stmt_3245/XOR_u32_u32_3233_Sample/$exit
      -- 	branch_block_stmt_2042/assign_stmt_3175_to_assign_stmt_3245/XOR_u32_u32_3233_Sample/ra
      -- 
    ra_13611_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => XOR_u32_u32_3233_inst_ack_0, ack => cp_elements(794)); -- 
    -- CP-element group 795 transition  input  output  bypass 
    -- predecessors 791 
    -- successors 797 
    -- members (10) 
      -- 	branch_block_stmt_2042/assign_stmt_3175_to_assign_stmt_3245/XOR_u32_u32_3233_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3175_to_assign_stmt_3245/XOR_u32_u32_3233_Update/$exit
      -- 	branch_block_stmt_2042/assign_stmt_3175_to_assign_stmt_3245/XOR_u32_u32_3233_Update/ca
      -- 	branch_block_stmt_2042/assign_stmt_3175_to_assign_stmt_3245/AND_u32_u32_3239_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_3175_to_assign_stmt_3245/R_iNsTr_98_3236_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_3175_to_assign_stmt_3245/R_iNsTr_98_3236_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3175_to_assign_stmt_3245/R_iNsTr_98_3236_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_3175_to_assign_stmt_3245/R_iNsTr_98_3236_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3175_to_assign_stmt_3245/AND_u32_u32_3239_Sample/$entry
      -- 	branch_block_stmt_2042/assign_stmt_3175_to_assign_stmt_3245/AND_u32_u32_3239_Sample/rr
      -- 
    ca_13616_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => XOR_u32_u32_3233_inst_ack_1, ack => cp_elements(795)); -- 
    rr_13628_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(795), ack => AND_u32_u32_3239_inst_req_0); -- 
    -- CP-element group 796 transition  output  bypass 
    -- predecessors 755 
    -- successors 798 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_3175_to_assign_stmt_3245/AND_u32_u32_3239_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_3175_to_assign_stmt_3245/AND_u32_u32_3239_Update/$entry
      -- 	branch_block_stmt_2042/assign_stmt_3175_to_assign_stmt_3245/AND_u32_u32_3239_Update/cr
      -- 
    cp_elements(796) <= cp_elements(755);
    cr_13633_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(796), ack => AND_u32_u32_3239_inst_req_1); -- 
    -- CP-element group 797 transition  input  bypass 
    -- predecessors 795 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_3175_to_assign_stmt_3245/AND_u32_u32_3239_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3175_to_assign_stmt_3245/AND_u32_u32_3239_Sample/$exit
      -- 	branch_block_stmt_2042/assign_stmt_3175_to_assign_stmt_3245/AND_u32_u32_3239_Sample/ra
      -- 
    ra_13629_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => AND_u32_u32_3239_inst_ack_0, ack => cp_elements(797)); -- 
    -- CP-element group 798 transition  input  bypass 
    -- predecessors 796 
    -- successors 803 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_3175_to_assign_stmt_3245/AND_u32_u32_3239_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3175_to_assign_stmt_3245/AND_u32_u32_3239_Update/$exit
      -- 	branch_block_stmt_2042/assign_stmt_3175_to_assign_stmt_3245/AND_u32_u32_3239_Update/ca
      -- 
    ca_13634_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => AND_u32_u32_3239_inst_ack_1, ack => cp_elements(798)); -- 
    -- CP-element group 799 join  transition  output  bypass 
    -- predecessors 762 769 
    -- successors 801 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_3175_to_assign_stmt_3245/SUB_u32_u32_3244_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_3175_to_assign_stmt_3245/SUB_u32_u32_3244_Sample/$entry
      -- 	branch_block_stmt_2042/assign_stmt_3175_to_assign_stmt_3245/SUB_u32_u32_3244_Sample/rr
      -- 
    cp_element_group_799: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 20) := "cp_element_group_799"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(762) & cp_elements(769);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(799), clk => clk, reset => reset); --
    end block;
    rr_13650_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(799), ack => SUB_u32_u32_3244_inst_req_0); -- 
    -- CP-element group 800 transition  output  bypass 
    -- predecessors 755 
    -- successors 802 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_3175_to_assign_stmt_3245/SUB_u32_u32_3244_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_3175_to_assign_stmt_3245/SUB_u32_u32_3244_Update/$entry
      -- 	branch_block_stmt_2042/assign_stmt_3175_to_assign_stmt_3245/SUB_u32_u32_3244_Update/cr
      -- 
    cp_elements(800) <= cp_elements(755);
    cr_13655_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(800), ack => SUB_u32_u32_3244_inst_req_1); -- 
    -- CP-element group 801 transition  input  bypass 
    -- predecessors 799 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_3175_to_assign_stmt_3245/SUB_u32_u32_3244_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3175_to_assign_stmt_3245/SUB_u32_u32_3244_Sample/$exit
      -- 	branch_block_stmt_2042/assign_stmt_3175_to_assign_stmt_3245/SUB_u32_u32_3244_Sample/ra
      -- 
    ra_13651_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => SUB_u32_u32_3244_inst_ack_0, ack => cp_elements(801)); -- 
    -- CP-element group 802 transition  input  bypass 
    -- predecessors 800 
    -- successors 803 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_3175_to_assign_stmt_3245/SUB_u32_u32_3244_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3175_to_assign_stmt_3245/SUB_u32_u32_3244_Update/$exit
      -- 	branch_block_stmt_2042/assign_stmt_3175_to_assign_stmt_3245/SUB_u32_u32_3244_Update/ca
      -- 
    ca_13656_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => SUB_u32_u32_3244_inst_ack_1, ack => cp_elements(802)); -- 
    -- CP-element group 803 join  transition  bypass 
    -- predecessors 779 789 798 802 
    -- successors 45 
    -- members (1) 
      -- 	branch_block_stmt_2042/assign_stmt_3175_to_assign_stmt_3245/$exit
      -- 
    cp_element_group_803: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 20) := "cp_element_group_803"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= cp_elements(779) & cp_elements(789) & cp_elements(798) & cp_elements(802);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(803), clk => clk, reset => reset); --
    end block;
    -- CP-element group 804 transition  place  dead  bypass 
    -- predecessors 45 
    -- successors 46 
    -- members (8) 
      -- 	branch_block_stmt_2042/merge_stmt_3256__entry__
      -- 	branch_block_stmt_2042/switch_stmt_3246__exit__
      -- 	branch_block_stmt_2042/switch_stmt_3246_dead_link/$entry
      -- 	branch_block_stmt_2042/switch_stmt_3246_dead_link/$exit
      -- 	branch_block_stmt_2042/switch_stmt_3246_dead_link/dead_transition
      -- 	branch_block_stmt_2042/merge_stmt_3256_dead_link/$entry
      -- 	branch_block_stmt_2042/merge_stmt_3256_dead_link/$exit
      -- 	branch_block_stmt_2042/merge_stmt_3256_dead_link/dead_transition
      -- 
    cp_elements(804) <= false;
    -- CP-element group 805 place  bypass 
    -- predecessors 45 
    -- successors 806 
    -- members (1) 
      -- 	branch_block_stmt_2042/switch_stmt_3246__condition_check_place__
      -- 
    cp_elements(805) <= cp_elements(45);
    -- CP-element group 806 fork  transition  bypass 
    -- predecessors 805 
    -- successors 807 813 
    -- members (1) 
      -- 	branch_block_stmt_2042/switch_stmt_3246__condition_check__/$entry
      -- 
    cp_elements(806) <= cp_elements(805);
    -- CP-element group 807 fork  transition  bypass 
    -- predecessors 806 
    -- successors 808 810 
    -- members (2) 
      -- 	branch_block_stmt_2042/switch_stmt_3246__condition_check__/condition_0/$entry
      -- 	branch_block_stmt_2042/switch_stmt_3246__condition_check__/condition_0/SplitProtocol/$entry
      -- 
    cp_elements(807) <= cp_elements(806);
    -- CP-element group 808 transition  output  bypass 
    -- predecessors 807 
    -- successors 809 
    -- members (2) 
      -- 	branch_block_stmt_2042/switch_stmt_3246__condition_check__/condition_0/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_2042/switch_stmt_3246__condition_check__/condition_0/SplitProtocol/Sample/rr
      -- 
    cp_elements(808) <= cp_elements(807);
    rr_13674_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(808), ack => switch_stmt_3246_select_expr_0_req_0); -- 
    -- CP-element group 809 transition  input  bypass 
    -- predecessors 808 
    -- successors 812 
    -- members (2) 
      -- 	branch_block_stmt_2042/switch_stmt_3246__condition_check__/condition_0/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_2042/switch_stmt_3246__condition_check__/condition_0/SplitProtocol/Sample/ra
      -- 
    ra_13675_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => switch_stmt_3246_select_expr_0_ack_0, ack => cp_elements(809)); -- 
    -- CP-element group 810 transition  output  bypass 
    -- predecessors 807 
    -- successors 811 
    -- members (2) 
      -- 	branch_block_stmt_2042/switch_stmt_3246__condition_check__/condition_0/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_2042/switch_stmt_3246__condition_check__/condition_0/SplitProtocol/Update/cr
      -- 
    cp_elements(810) <= cp_elements(807);
    cr_13679_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(810), ack => switch_stmt_3246_select_expr_0_req_1); -- 
    -- CP-element group 811 transition  input  bypass 
    -- predecessors 810 
    -- successors 812 
    -- members (2) 
      -- 	branch_block_stmt_2042/switch_stmt_3246__condition_check__/condition_0/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_2042/switch_stmt_3246__condition_check__/condition_0/SplitProtocol/Update/ca
      -- 
    ca_13680_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => switch_stmt_3246_select_expr_0_ack_1, ack => cp_elements(811)); -- 
    -- CP-element group 812 join  transition  output  bypass 
    -- predecessors 809 811 
    -- successors 819 
    -- members (3) 
      -- 	branch_block_stmt_2042/switch_stmt_3246__condition_check__/condition_0/$exit
      -- 	branch_block_stmt_2042/switch_stmt_3246__condition_check__/condition_0/SplitProtocol/$exit
      -- 	branch_block_stmt_2042/switch_stmt_3246__condition_check__/condition_0/cmp
      -- 
    cp_element_group_812: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 20) := "cp_element_group_812"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(809) & cp_elements(811);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(812), clk => clk, reset => reset); --
    end block;
    cmp_13681_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(812), ack => switch_stmt_3246_branch_0_req_0); -- 
    -- CP-element group 813 fork  transition  bypass 
    -- predecessors 806 
    -- successors 814 816 
    -- members (2) 
      -- 	branch_block_stmt_2042/switch_stmt_3246__condition_check__/condition_1/$entry
      -- 	branch_block_stmt_2042/switch_stmt_3246__condition_check__/condition_1/SplitProtocol/$entry
      -- 
    cp_elements(813) <= cp_elements(806);
    -- CP-element group 814 transition  output  bypass 
    -- predecessors 813 
    -- successors 815 
    -- members (2) 
      -- 	branch_block_stmt_2042/switch_stmt_3246__condition_check__/condition_1/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_2042/switch_stmt_3246__condition_check__/condition_1/SplitProtocol/Sample/rr
      -- 
    cp_elements(814) <= cp_elements(813);
    rr_13691_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(814), ack => switch_stmt_3246_select_expr_1_req_0); -- 
    -- CP-element group 815 transition  input  bypass 
    -- predecessors 814 
    -- successors 818 
    -- members (2) 
      -- 	branch_block_stmt_2042/switch_stmt_3246__condition_check__/condition_1/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_2042/switch_stmt_3246__condition_check__/condition_1/SplitProtocol/Sample/ra
      -- 
    ra_13692_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => switch_stmt_3246_select_expr_1_ack_0, ack => cp_elements(815)); -- 
    -- CP-element group 816 transition  output  bypass 
    -- predecessors 813 
    -- successors 817 
    -- members (2) 
      -- 	branch_block_stmt_2042/switch_stmt_3246__condition_check__/condition_1/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_2042/switch_stmt_3246__condition_check__/condition_1/SplitProtocol/Update/cr
      -- 
    cp_elements(816) <= cp_elements(813);
    cr_13696_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(816), ack => switch_stmt_3246_select_expr_1_req_1); -- 
    -- CP-element group 817 transition  input  bypass 
    -- predecessors 816 
    -- successors 818 
    -- members (2) 
      -- 	branch_block_stmt_2042/switch_stmt_3246__condition_check__/condition_1/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_2042/switch_stmt_3246__condition_check__/condition_1/SplitProtocol/Update/ca
      -- 
    ca_13697_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => switch_stmt_3246_select_expr_1_ack_1, ack => cp_elements(817)); -- 
    -- CP-element group 818 join  transition  output  bypass 
    -- predecessors 815 817 
    -- successors 819 
    -- members (3) 
      -- 	branch_block_stmt_2042/switch_stmt_3246__condition_check__/condition_1/$exit
      -- 	branch_block_stmt_2042/switch_stmt_3246__condition_check__/condition_1/SplitProtocol/$exit
      -- 	branch_block_stmt_2042/switch_stmt_3246__condition_check__/condition_1/cmp
      -- 
    cp_element_group_818: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 20) := "cp_element_group_818"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(815) & cp_elements(817);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(818), clk => clk, reset => reset); --
    end block;
    cmp_13698_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(818), ack => switch_stmt_3246_branch_1_req_0); -- 
    -- CP-element group 819 join  transition  output  bypass 
    -- predecessors 812 818 
    -- successors 820 
    -- members (1) 
      -- 	branch_block_stmt_2042/switch_stmt_3246__condition_check__/$exit
      -- 
    cp_element_group_819: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 20) := "cp_element_group_819"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(812) & cp_elements(818);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(819), clk => clk, reset => reset); --
    end block;
    Xexit_13664_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(819), ack => switch_stmt_3246_branch_default_req_0); -- 
    -- CP-element group 820 branch  place  bypass 
    -- predecessors 819 
    -- successors 821 823 825 
    -- members (1) 
      -- 	branch_block_stmt_2042/switch_stmt_3246__select__
      -- 
    cp_elements(820) <= cp_elements(819);
    -- CP-element group 821 transition  bypass 
    -- predecessors 820 
    -- successors 822 
    -- members (1) 
      -- 	branch_block_stmt_2042/switch_stmt_3246_choice_0/$entry
      -- 
    cp_elements(821) <= cp_elements(820);
    -- CP-element group 822 fork  transition  place  input  bypass 
    -- predecessors 821 
    -- successors 2136 2137 
    -- members (8) 
      -- 	branch_block_stmt_2042/switch_stmt_3246_choice_0/$exit
      -- 	branch_block_stmt_2042/switch_stmt_3246_choice_0/ack1
      -- 	branch_block_stmt_2042/bb_41_xx_xloopexitx_xix_xix_xi
      -- 	branch_block_stmt_2042/bb_41_xx_xloopexitx_xix_xix_xi_PhiReq/$entry
      -- 	branch_block_stmt_2042/bb_41_xx_xloopexitx_xix_xix_xi_PhiReq/phi_stmt_3385/$entry
      -- 	branch_block_stmt_2042/bb_41_xx_xloopexitx_xix_xix_xi_PhiReq/phi_stmt_3385/phi_stmt_3385_sources/$entry
      -- 	branch_block_stmt_2042/bb_41_xx_xloopexitx_xix_xix_xi_PhiReq/phi_stmt_3385/phi_stmt_3385_sources/type_cast_3391/$entry
      -- 	branch_block_stmt_2042/bb_41_xx_xloopexitx_xix_xix_xi_PhiReq/phi_stmt_3385/phi_stmt_3385_sources/type_cast_3391/SplitProtocol/$entry
      -- 
    ack1_13703_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => switch_stmt_3246_branch_0_ack_1, ack => cp_elements(822)); -- 
    -- CP-element group 823 transition  bypass 
    -- predecessors 820 
    -- successors 824 
    -- members (1) 
      -- 	branch_block_stmt_2042/switch_stmt_3246_choice_1/$entry
      -- 
    cp_elements(823) <= cp_elements(820);
    -- CP-element group 824 fork  transition  place  input  bypass 
    -- predecessors 823 
    -- successors 2147 2151 
    -- members (6) 
      -- 	branch_block_stmt_2042/switch_stmt_3246_choice_1/$exit
      -- 	branch_block_stmt_2042/switch_stmt_3246_choice_1/ack1
      -- 	branch_block_stmt_2042/bb_41_udiv32x_xexitx_xpreheaderx_xix_xi
      -- 	branch_block_stmt_2042/bb_41_udiv32x_xexitx_xpreheaderx_xix_xi_PhiReq/phi_stmt_3395/phi_stmt_3395_sources/$entry
      -- 	branch_block_stmt_2042/bb_41_udiv32x_xexitx_xpreheaderx_xix_xi_PhiReq/phi_stmt_3395/$entry
      -- 	branch_block_stmt_2042/bb_41_udiv32x_xexitx_xpreheaderx_xix_xi_PhiReq/$entry
      -- 
    ack1_13708_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => switch_stmt_3246_branch_1_ack_1, ack => cp_elements(824)); -- 
    -- CP-element group 825 transition  bypass 
    -- predecessors 820 
    -- successors 826 
    -- members (1) 
      -- 	branch_block_stmt_2042/switch_stmt_3246_choice_default/$entry
      -- 
    cp_elements(825) <= cp_elements(820);
    -- CP-element group 826 transition  place  input  bypass 
    -- predecessors 825 
    -- successors 46 
    -- members (9) 
      -- 	branch_block_stmt_2042/switch_stmt_3246_choice_default/$exit
      -- 	branch_block_stmt_2042/switch_stmt_3246_choice_default/ack0
      -- 	branch_block_stmt_2042/bb_41_bbx_xnph7x_xix_xix_xix_xpreheader
      -- 	branch_block_stmt_2042/merge_stmt_3256_PhiReqMerge
      -- 	branch_block_stmt_2042/bb_41_bbx_xnph7x_xix_xix_xix_xpreheader_PhiReq/$entry
      -- 	branch_block_stmt_2042/bb_41_bbx_xnph7x_xix_xix_xix_xpreheader_PhiReq/$exit
      -- 	branch_block_stmt_2042/merge_stmt_3256_PhiAck/$entry
      -- 	branch_block_stmt_2042/merge_stmt_3256_PhiAck/$exit
      -- 	branch_block_stmt_2042/merge_stmt_3256_PhiAck/dummy
      -- 
    ack0_13713_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => switch_stmt_3246_branch_default_ack_0, ack => cp_elements(826)); -- 
    -- CP-element group 827 fork  transition  bypass 
    -- predecessors 47 
    -- successors 828 829 833 834 
    -- members (1) 
      -- 	branch_block_stmt_2042/assign_stmt_3278_to_assign_stmt_3283/$entry
      -- 
    cp_elements(827) <= cp_elements(47);
    -- CP-element group 828 transition  output  bypass 
    -- predecessors 827 
    -- successors 831 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_3278_to_assign_stmt_3283/LSHR_u32_u32_3277_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_3278_to_assign_stmt_3283/LSHR_u32_u32_3277_Update/$entry
      -- 	branch_block_stmt_2042/assign_stmt_3278_to_assign_stmt_3283/LSHR_u32_u32_3277_Update/cr
      -- 
    cp_elements(828) <= cp_elements(827);
    cr_13734_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(828), ack => LSHR_u32_u32_3277_inst_req_1); -- 
    -- CP-element group 829 transition  output  bypass 
    -- predecessors 827 
    -- successors 830 
    -- members (7) 
      -- 	branch_block_stmt_2042/assign_stmt_3278_to_assign_stmt_3283/LSHR_u32_u32_3277_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_3278_to_assign_stmt_3283/R_xx_x016x_xix_xix_xi_3274_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_3278_to_assign_stmt_3283/R_xx_x016x_xix_xix_xi_3274_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3278_to_assign_stmt_3283/R_xx_x016x_xix_xix_xi_3274_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_3278_to_assign_stmt_3283/R_xx_x016x_xix_xix_xi_3274_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3278_to_assign_stmt_3283/LSHR_u32_u32_3277_Sample/$entry
      -- 	branch_block_stmt_2042/assign_stmt_3278_to_assign_stmt_3283/LSHR_u32_u32_3277_Sample/rr
      -- 
    cp_elements(829) <= cp_elements(827);
    rr_13729_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(829), ack => LSHR_u32_u32_3277_inst_req_0); -- 
    -- CP-element group 830 transition  input  bypass 
    -- predecessors 829 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_3278_to_assign_stmt_3283/LSHR_u32_u32_3277_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3278_to_assign_stmt_3283/LSHR_u32_u32_3277_Sample/$exit
      -- 	branch_block_stmt_2042/assign_stmt_3278_to_assign_stmt_3283/LSHR_u32_u32_3277_Sample/ra
      -- 
    ra_13730_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => LSHR_u32_u32_3277_inst_ack_0, ack => cp_elements(830)); -- 
    -- CP-element group 831 transition  input  bypass 
    -- predecessors 828 
    -- successors 832 
    -- members (7) 
      -- 	branch_block_stmt_2042/assign_stmt_3278_to_assign_stmt_3283/LSHR_u32_u32_3277_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3278_to_assign_stmt_3283/LSHR_u32_u32_3277_Update/$exit
      -- 	branch_block_stmt_2042/assign_stmt_3278_to_assign_stmt_3283/LSHR_u32_u32_3277_Update/ca
      -- 	branch_block_stmt_2042/assign_stmt_3278_to_assign_stmt_3283/R_iNsTr_154_3280_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_3278_to_assign_stmt_3283/R_iNsTr_154_3280_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3278_to_assign_stmt_3283/R_iNsTr_154_3280_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_3278_to_assign_stmt_3283/R_iNsTr_154_3280_update_completed_
      -- 
    ca_13735_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => LSHR_u32_u32_3277_inst_ack_1, ack => cp_elements(831)); -- 
    -- CP-element group 832 join  transition  output  bypass 
    -- predecessors 831 834 
    -- successors 835 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_3278_to_assign_stmt_3283/UGT_u32_u1_3282_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_3278_to_assign_stmt_3283/UGT_u32_u1_3282_Sample/$entry
      -- 	branch_block_stmt_2042/assign_stmt_3278_to_assign_stmt_3283/UGT_u32_u1_3282_Sample/rr
      -- 
    cp_element_group_832: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 20) := "cp_element_group_832"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(831) & cp_elements(834);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(832), clk => clk, reset => reset); --
    end block;
    rr_13751_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(832), ack => UGT_u32_u1_3282_inst_req_0); -- 
    -- CP-element group 833 transition  output  bypass 
    -- predecessors 827 
    -- successors 836 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_3278_to_assign_stmt_3283/UGT_u32_u1_3282_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_3278_to_assign_stmt_3283/UGT_u32_u1_3282_Update/$entry
      -- 	branch_block_stmt_2042/assign_stmt_3278_to_assign_stmt_3283/UGT_u32_u1_3282_Update/cr
      -- 
    cp_elements(833) <= cp_elements(827);
    cr_13756_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(833), ack => UGT_u32_u1_3282_inst_req_1); -- 
    -- CP-element group 834 transition  bypass 
    -- predecessors 827 
    -- successors 832 
    -- members (4) 
      -- 	branch_block_stmt_2042/assign_stmt_3278_to_assign_stmt_3283/R_iNsTr_97_3281_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_3278_to_assign_stmt_3283/R_iNsTr_97_3281_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3278_to_assign_stmt_3283/R_iNsTr_97_3281_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_3278_to_assign_stmt_3283/R_iNsTr_97_3281_update_completed_
      -- 
    cp_elements(834) <= cp_elements(827);
    -- CP-element group 835 transition  input  bypass 
    -- predecessors 832 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_3278_to_assign_stmt_3283/UGT_u32_u1_3282_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3278_to_assign_stmt_3283/UGT_u32_u1_3282_Sample/$exit
      -- 	branch_block_stmt_2042/assign_stmt_3278_to_assign_stmt_3283/UGT_u32_u1_3282_Sample/ra
      -- 
    ra_13752_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => UGT_u32_u1_3282_inst_ack_0, ack => cp_elements(835)); -- 
    -- CP-element group 836 branch  transition  place  input  bypass 
    -- predecessors 833 
    -- successors 837 838 
    -- members (6) 
      -- 	branch_block_stmt_2042/assign_stmt_3278_to_assign_stmt_3283__exit__
      -- 	branch_block_stmt_2042/if_stmt_3284__entry__
      -- 	branch_block_stmt_2042/assign_stmt_3278_to_assign_stmt_3283/$exit
      -- 	branch_block_stmt_2042/assign_stmt_3278_to_assign_stmt_3283/UGT_u32_u1_3282_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3278_to_assign_stmt_3283/UGT_u32_u1_3282_Update/$exit
      -- 	branch_block_stmt_2042/assign_stmt_3278_to_assign_stmt_3283/UGT_u32_u1_3282_Update/ca
      -- 
    ca_13757_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => UGT_u32_u1_3282_inst_ack_1, ack => cp_elements(836)); -- 
    -- CP-element group 837 transition  place  dead  bypass 
    -- predecessors 836 
    -- successors 48 
    -- members (8) 
      -- 	branch_block_stmt_2042/if_stmt_3284__exit__
      -- 	branch_block_stmt_2042/merge_stmt_3290__entry__
      -- 	branch_block_stmt_2042/if_stmt_3284_dead_link/$entry
      -- 	branch_block_stmt_2042/if_stmt_3284_dead_link/$exit
      -- 	branch_block_stmt_2042/if_stmt_3284_dead_link/dead_transition
      -- 	branch_block_stmt_2042/merge_stmt_3290_dead_link/$entry
      -- 	branch_block_stmt_2042/merge_stmt_3290_dead_link/$exit
      -- 	branch_block_stmt_2042/merge_stmt_3290_dead_link/dead_transition
      -- 
    cp_elements(837) <= false;
    -- CP-element group 838 transition  output  bypass 
    -- predecessors 836 
    -- successors 839 
    -- members (3) 
      -- 	branch_block_stmt_2042/if_stmt_3284_eval_test/$entry
      -- 	branch_block_stmt_2042/if_stmt_3284_eval_test/$exit
      -- 	branch_block_stmt_2042/if_stmt_3284_eval_test/branch_req
      -- 
    cp_elements(838) <= cp_elements(836);
    branch_req_13765_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(838), ack => if_stmt_3284_branch_req_0); -- 
    -- CP-element group 839 branch  place  bypass 
    -- predecessors 838 
    -- successors 840 842 
    -- members (1) 
      -- 	branch_block_stmt_2042/R_iNsTr_155_3285_place
      -- 
    cp_elements(839) <= cp_elements(838);
    -- CP-element group 840 transition  bypass 
    -- predecessors 839 
    -- successors 841 
    -- members (1) 
      -- 	branch_block_stmt_2042/if_stmt_3284_if_link/$entry
      -- 
    cp_elements(840) <= cp_elements(839);
    -- CP-element group 841 transition  place  input  bypass 
    -- predecessors 840 
    -- successors 48 
    -- members (9) 
      -- 	branch_block_stmt_2042/if_stmt_3284_if_link/$exit
      -- 	branch_block_stmt_2042/if_stmt_3284_if_link/if_choice_transition
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xix_xi_bbx_xnphx_xix_xix_xix_xpreheader
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xix_xi_bbx_xnphx_xix_xix_xix_xpreheader_PhiReq/$entry
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xix_xi_bbx_xnphx_xix_xix_xix_xpreheader_PhiReq/$exit
      -- 	branch_block_stmt_2042/merge_stmt_3290_PhiReqMerge
      -- 	branch_block_stmt_2042/merge_stmt_3290_PhiAck/$entry
      -- 	branch_block_stmt_2042/merge_stmt_3290_PhiAck/$exit
      -- 	branch_block_stmt_2042/merge_stmt_3290_PhiAck/dummy
      -- 
    if_choice_transition_13770_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_3284_branch_ack_1, ack => cp_elements(841)); -- 
    -- CP-element group 842 transition  bypass 
    -- predecessors 839 
    -- successors 843 
    -- members (1) 
      -- 	branch_block_stmt_2042/if_stmt_3284_else_link/$entry
      -- 
    cp_elements(842) <= cp_elements(839);
    -- CP-element group 843 transition  place  input  bypass 
    -- predecessors 842 
    -- successors 2087 
    -- members (3) 
      -- 	branch_block_stmt_2042/if_stmt_3284_else_link/$exit
      -- 	branch_block_stmt_2042/if_stmt_3284_else_link/else_choice_transition
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xix_xi_xx_x_crit_edgex_xix_xix_xi
      -- 
    else_choice_transition_13774_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_3284_branch_ack_0, ack => cp_elements(843)); -- 
    -- CP-element group 844 fork  transition  bypass 
    -- predecessors 49 
    -- successors 845 846 849 850 854 855 
    -- members (1) 
      -- 	branch_block_stmt_2042/assign_stmt_3312_to_assign_stmt_3323/$entry
      -- 
    cp_elements(844) <= cp_elements(49);
    -- CP-element group 845 transition  output  bypass 
    -- predecessors 844 
    -- successors 848 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_3312_to_assign_stmt_3323/SHL_u32_u32_3311_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_3312_to_assign_stmt_3323/SHL_u32_u32_3311_Update/$entry
      -- 	branch_block_stmt_2042/assign_stmt_3312_to_assign_stmt_3323/SHL_u32_u32_3311_Update/cr
      -- 
    cp_elements(845) <= cp_elements(844);
    cr_13796_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(845), ack => SHL_u32_u32_3311_inst_req_1); -- 
    -- CP-element group 846 transition  output  bypass 
    -- predecessors 844 
    -- successors 847 
    -- members (7) 
      -- 	branch_block_stmt_2042/assign_stmt_3312_to_assign_stmt_3323/SHL_u32_u32_3311_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_3312_to_assign_stmt_3323/R_shifted_divisorx_x03x_xix_xix_xi_3308_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_3312_to_assign_stmt_3323/R_shifted_divisorx_x03x_xix_xix_xi_3308_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3312_to_assign_stmt_3323/R_shifted_divisorx_x03x_xix_xix_xi_3308_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_3312_to_assign_stmt_3323/R_shifted_divisorx_x03x_xix_xix_xi_3308_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3312_to_assign_stmt_3323/SHL_u32_u32_3311_Sample/$entry
      -- 	branch_block_stmt_2042/assign_stmt_3312_to_assign_stmt_3323/SHL_u32_u32_3311_Sample/rr
      -- 
    cp_elements(846) <= cp_elements(844);
    rr_13791_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(846), ack => SHL_u32_u32_3311_inst_req_0); -- 
    -- CP-element group 847 transition  input  bypass 
    -- predecessors 846 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_3312_to_assign_stmt_3323/SHL_u32_u32_3311_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3312_to_assign_stmt_3323/SHL_u32_u32_3311_Sample/$exit
      -- 	branch_block_stmt_2042/assign_stmt_3312_to_assign_stmt_3323/SHL_u32_u32_3311_Sample/ra
      -- 
    ra_13792_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => SHL_u32_u32_3311_inst_ack_0, ack => cp_elements(847)); -- 
    -- CP-element group 848 transition  input  bypass 
    -- predecessors 845 
    -- successors 853 
    -- members (7) 
      -- 	branch_block_stmt_2042/assign_stmt_3312_to_assign_stmt_3323/SHL_u32_u32_3311_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3312_to_assign_stmt_3323/SHL_u32_u32_3311_Update/$exit
      -- 	branch_block_stmt_2042/assign_stmt_3312_to_assign_stmt_3323/SHL_u32_u32_3311_Update/ca
      -- 	branch_block_stmt_2042/assign_stmt_3312_to_assign_stmt_3323/R_iNsTr_226_3320_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_3312_to_assign_stmt_3323/R_iNsTr_226_3320_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3312_to_assign_stmt_3323/R_iNsTr_226_3320_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_3312_to_assign_stmt_3323/R_iNsTr_226_3320_update_completed_
      -- 
    ca_13797_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => SHL_u32_u32_3311_inst_ack_1, ack => cp_elements(848)); -- 
    -- CP-element group 849 transition  output  bypass 
    -- predecessors 844 
    -- successors 852 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_3312_to_assign_stmt_3323/SHL_u32_u32_3317_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_3312_to_assign_stmt_3323/SHL_u32_u32_3317_Update/$entry
      -- 	branch_block_stmt_2042/assign_stmt_3312_to_assign_stmt_3323/SHL_u32_u32_3317_Update/cr
      -- 
    cp_elements(849) <= cp_elements(844);
    cr_13814_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(849), ack => SHL_u32_u32_3317_inst_req_1); -- 
    -- CP-element group 850 transition  output  bypass 
    -- predecessors 844 
    -- successors 851 
    -- members (7) 
      -- 	branch_block_stmt_2042/assign_stmt_3312_to_assign_stmt_3323/SHL_u32_u32_3317_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_3312_to_assign_stmt_3323/R_curr_quotientx_x02x_xix_xix_xi_3314_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_3312_to_assign_stmt_3323/R_curr_quotientx_x02x_xix_xix_xi_3314_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3312_to_assign_stmt_3323/R_curr_quotientx_x02x_xix_xix_xi_3314_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_3312_to_assign_stmt_3323/R_curr_quotientx_x02x_xix_xix_xi_3314_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3312_to_assign_stmt_3323/SHL_u32_u32_3317_Sample/$entry
      -- 	branch_block_stmt_2042/assign_stmt_3312_to_assign_stmt_3323/SHL_u32_u32_3317_Sample/rr
      -- 
    cp_elements(850) <= cp_elements(844);
    rr_13809_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(850), ack => SHL_u32_u32_3317_inst_req_0); -- 
    -- CP-element group 851 transition  input  bypass 
    -- predecessors 850 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_3312_to_assign_stmt_3323/SHL_u32_u32_3317_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3312_to_assign_stmt_3323/SHL_u32_u32_3317_Sample/$exit
      -- 	branch_block_stmt_2042/assign_stmt_3312_to_assign_stmt_3323/SHL_u32_u32_3317_Sample/ra
      -- 
    ra_13810_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => SHL_u32_u32_3317_inst_ack_0, ack => cp_elements(851)); -- 
    -- CP-element group 852 transition  input  bypass 
    -- predecessors 849 
    -- successors 858 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_3312_to_assign_stmt_3323/SHL_u32_u32_3317_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3312_to_assign_stmt_3323/SHL_u32_u32_3317_Update/$exit
      -- 	branch_block_stmt_2042/assign_stmt_3312_to_assign_stmt_3323/SHL_u32_u32_3317_Update/ca
      -- 
    ca_13815_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => SHL_u32_u32_3317_inst_ack_1, ack => cp_elements(852)); -- 
    -- CP-element group 853 join  transition  output  bypass 
    -- predecessors 848 855 
    -- successors 856 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_3312_to_assign_stmt_3323/ULT_u32_u1_3322_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_3312_to_assign_stmt_3323/ULT_u32_u1_3322_Sample/$entry
      -- 	branch_block_stmt_2042/assign_stmt_3312_to_assign_stmt_3323/ULT_u32_u1_3322_Sample/rr
      -- 
    cp_element_group_853: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 20) := "cp_element_group_853"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(848) & cp_elements(855);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(853), clk => clk, reset => reset); --
    end block;
    rr_13831_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(853), ack => ULT_u32_u1_3322_inst_req_0); -- 
    -- CP-element group 854 transition  output  bypass 
    -- predecessors 844 
    -- successors 857 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_3312_to_assign_stmt_3323/ULT_u32_u1_3322_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_3312_to_assign_stmt_3323/ULT_u32_u1_3322_Update/$entry
      -- 	branch_block_stmt_2042/assign_stmt_3312_to_assign_stmt_3323/ULT_u32_u1_3322_Update/cr
      -- 
    cp_elements(854) <= cp_elements(844);
    cr_13836_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(854), ack => ULT_u32_u1_3322_inst_req_1); -- 
    -- CP-element group 855 transition  bypass 
    -- predecessors 844 
    -- successors 853 
    -- members (4) 
      -- 	branch_block_stmt_2042/assign_stmt_3312_to_assign_stmt_3323/R_iNsTr_154_3321_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_3312_to_assign_stmt_3323/R_iNsTr_154_3321_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3312_to_assign_stmt_3323/R_iNsTr_154_3321_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_3312_to_assign_stmt_3323/R_iNsTr_154_3321_update_completed_
      -- 
    cp_elements(855) <= cp_elements(844);
    -- CP-element group 856 transition  input  bypass 
    -- predecessors 853 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_3312_to_assign_stmt_3323/ULT_u32_u1_3322_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3312_to_assign_stmt_3323/ULT_u32_u1_3322_Sample/$exit
      -- 	branch_block_stmt_2042/assign_stmt_3312_to_assign_stmt_3323/ULT_u32_u1_3322_Sample/ra
      -- 
    ra_13832_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ULT_u32_u1_3322_inst_ack_0, ack => cp_elements(856)); -- 
    -- CP-element group 857 transition  input  bypass 
    -- predecessors 854 
    -- successors 858 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_3312_to_assign_stmt_3323/ULT_u32_u1_3322_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3312_to_assign_stmt_3323/ULT_u32_u1_3322_Update/$exit
      -- 	branch_block_stmt_2042/assign_stmt_3312_to_assign_stmt_3323/ULT_u32_u1_3322_Update/ca
      -- 
    ca_13837_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ULT_u32_u1_3322_inst_ack_1, ack => cp_elements(857)); -- 
    -- CP-element group 858 join  transition  bypass 
    -- predecessors 852 857 
    -- successors 50 
    -- members (1) 
      -- 	branch_block_stmt_2042/assign_stmt_3312_to_assign_stmt_3323/$exit
      -- 
    cp_element_group_858: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 20) := "cp_element_group_858"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(852) & cp_elements(857);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(858), clk => clk, reset => reset); --
    end block;
    -- CP-element group 859 transition  place  dead  bypass 
    -- predecessors 50 
    -- successors 51 
    -- members (8) 
      -- 	branch_block_stmt_2042/merge_stmt_3330__entry__
      -- 	branch_block_stmt_2042/if_stmt_3324__exit__
      -- 	branch_block_stmt_2042/if_stmt_3324_dead_link/$entry
      -- 	branch_block_stmt_2042/if_stmt_3324_dead_link/$exit
      -- 	branch_block_stmt_2042/if_stmt_3324_dead_link/dead_transition
      -- 	branch_block_stmt_2042/merge_stmt_3330_dead_link/$entry
      -- 	branch_block_stmt_2042/merge_stmt_3330_dead_link/$exit
      -- 	branch_block_stmt_2042/merge_stmt_3330_dead_link/dead_transition
      -- 
    cp_elements(859) <= false;
    -- CP-element group 860 transition  output  bypass 
    -- predecessors 50 
    -- successors 861 
    -- members (3) 
      -- 	branch_block_stmt_2042/if_stmt_3324_eval_test/$entry
      -- 	branch_block_stmt_2042/if_stmt_3324_eval_test/$exit
      -- 	branch_block_stmt_2042/if_stmt_3324_eval_test/branch_req
      -- 
    cp_elements(860) <= cp_elements(50);
    branch_req_13845_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(860), ack => if_stmt_3324_branch_req_0); -- 
    -- CP-element group 861 branch  place  bypass 
    -- predecessors 860 
    -- successors 862 864 
    -- members (1) 
      -- 	branch_block_stmt_2042/R_iNsTr_228_3325_place
      -- 
    cp_elements(861) <= cp_elements(860);
    -- CP-element group 862 transition  bypass 
    -- predecessors 861 
    -- successors 863 
    -- members (1) 
      -- 	branch_block_stmt_2042/if_stmt_3324_if_link/$entry
      -- 
    cp_elements(862) <= cp_elements(861);
    -- CP-element group 863 transition  place  input  bypass 
    -- predecessors 862 
    -- successors 2025 
    -- members (3) 
      -- 	branch_block_stmt_2042/if_stmt_3324_if_link/$exit
      -- 	branch_block_stmt_2042/if_stmt_3324_if_link/if_choice_transition
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi_bbx_xnphx_xix_xix_xi
      -- 
    if_choice_transition_13850_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_3324_branch_ack_1, ack => cp_elements(863)); -- 
    -- CP-element group 864 transition  bypass 
    -- predecessors 861 
    -- successors 865 
    -- members (1) 
      -- 	branch_block_stmt_2042/if_stmt_3324_else_link/$entry
      -- 
    cp_elements(864) <= cp_elements(861);
    -- CP-element group 865 transition  place  input  bypass 
    -- predecessors 864 
    -- successors 2068 
    -- members (3) 
      -- 	branch_block_stmt_2042/if_stmt_3324_else_link/$exit
      -- 	branch_block_stmt_2042/if_stmt_3324_else_link/else_choice_transition
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi_xx_x_crit_edgex_xix_xix_xix_xloopexit
      -- 
    else_choice_transition_13854_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_3324_branch_ack_0, ack => cp_elements(865)); -- 
    -- CP-element group 866 fork  transition  bypass 
    -- predecessors 52 
    -- successors 868 869 870 874 875 876 880 881 
    -- members (1) 
      -- 	branch_block_stmt_2042/assign_stmt_3360_to_assign_stmt_3370/$entry
      -- 
    cp_elements(866) <= cp_elements(52);
    -- CP-element group 867 join  transition  output  bypass 
    -- predecessors 869 870 
    -- successors 871 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_3360_to_assign_stmt_3370/ADD_u32_u32_3359_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_3360_to_assign_stmt_3370/ADD_u32_u32_3359_Sample/$entry
      -- 	branch_block_stmt_2042/assign_stmt_3360_to_assign_stmt_3370/ADD_u32_u32_3359_Sample/rr
      -- 
    cp_element_group_867: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 20) := "cp_element_group_867"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(869) & cp_elements(870);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(867), clk => clk, reset => reset); --
    end block;
    rr_13875_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(867), ack => ADD_u32_u32_3359_inst_req_0); -- 
    -- CP-element group 868 transition  output  bypass 
    -- predecessors 866 
    -- successors 872 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_3360_to_assign_stmt_3370/ADD_u32_u32_3359_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_3360_to_assign_stmt_3370/ADD_u32_u32_3359_Update/$entry
      -- 	branch_block_stmt_2042/assign_stmt_3360_to_assign_stmt_3370/ADD_u32_u32_3359_Update/cr
      -- 
    cp_elements(868) <= cp_elements(866);
    cr_13880_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(868), ack => ADD_u32_u32_3359_inst_req_1); -- 
    -- CP-element group 869 transition  bypass 
    -- predecessors 866 
    -- successors 867 
    -- members (4) 
      -- 	branch_block_stmt_2042/assign_stmt_3360_to_assign_stmt_3370/R_curr_quotientx_x0x_xlcssax_xix_xix_xi_3357_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_3360_to_assign_stmt_3370/R_curr_quotientx_x0x_xlcssax_xix_xix_xi_3357_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3360_to_assign_stmt_3370/R_curr_quotientx_x0x_xlcssax_xix_xix_xi_3357_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_3360_to_assign_stmt_3370/R_curr_quotientx_x0x_xlcssax_xix_xix_xi_3357_update_completed_
      -- 
    cp_elements(869) <= cp_elements(866);
    -- CP-element group 870 transition  bypass 
    -- predecessors 866 
    -- successors 867 
    -- members (4) 
      -- 	branch_block_stmt_2042/assign_stmt_3360_to_assign_stmt_3370/R_quotientx_x05x_xix_xix_xi_3358_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_3360_to_assign_stmt_3370/R_quotientx_x05x_xix_xix_xi_3358_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3360_to_assign_stmt_3370/R_quotientx_x05x_xix_xix_xi_3358_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_3360_to_assign_stmt_3370/R_quotientx_x05x_xix_xix_xi_3358_update_completed_
      -- 
    cp_elements(870) <= cp_elements(866);
    -- CP-element group 871 transition  input  bypass 
    -- predecessors 867 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_3360_to_assign_stmt_3370/ADD_u32_u32_3359_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3360_to_assign_stmt_3370/ADD_u32_u32_3359_Sample/$exit
      -- 	branch_block_stmt_2042/assign_stmt_3360_to_assign_stmt_3370/ADD_u32_u32_3359_Sample/ra
      -- 
    ra_13876_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u32_u32_3359_inst_ack_0, ack => cp_elements(871)); -- 
    -- CP-element group 872 transition  input  bypass 
    -- predecessors 868 
    -- successors 884 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_3360_to_assign_stmt_3370/ADD_u32_u32_3359_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3360_to_assign_stmt_3370/ADD_u32_u32_3359_Update/$exit
      -- 	branch_block_stmt_2042/assign_stmt_3360_to_assign_stmt_3370/ADD_u32_u32_3359_Update/ca
      -- 
    ca_13881_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u32_u32_3359_inst_ack_1, ack => cp_elements(872)); -- 
    -- CP-element group 873 join  transition  output  bypass 
    -- predecessors 875 876 
    -- successors 877 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_3360_to_assign_stmt_3370/SUB_u32_u32_3364_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_3360_to_assign_stmt_3370/SUB_u32_u32_3364_Sample/$entry
      -- 	branch_block_stmt_2042/assign_stmt_3360_to_assign_stmt_3370/SUB_u32_u32_3364_Sample/rr
      -- 
    cp_element_group_873: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 20) := "cp_element_group_873"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(875) & cp_elements(876);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(873), clk => clk, reset => reset); --
    end block;
    rr_13897_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(873), ack => SUB_u32_u32_3364_inst_req_0); -- 
    -- CP-element group 874 transition  output  bypass 
    -- predecessors 866 
    -- successors 878 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_3360_to_assign_stmt_3370/SUB_u32_u32_3364_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_3360_to_assign_stmt_3370/SUB_u32_u32_3364_Update/$entry
      -- 	branch_block_stmt_2042/assign_stmt_3360_to_assign_stmt_3370/SUB_u32_u32_3364_Update/cr
      -- 
    cp_elements(874) <= cp_elements(866);
    cr_13902_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(874), ack => SUB_u32_u32_3364_inst_req_1); -- 
    -- CP-element group 875 transition  bypass 
    -- predecessors 866 
    -- successors 873 
    -- members (4) 
      -- 	branch_block_stmt_2042/assign_stmt_3360_to_assign_stmt_3370/R_xx_x016x_xix_xix_xi_3362_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_3360_to_assign_stmt_3370/R_xx_x016x_xix_xix_xi_3362_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3360_to_assign_stmt_3370/R_xx_x016x_xix_xix_xi_3362_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_3360_to_assign_stmt_3370/R_xx_x016x_xix_xix_xi_3362_update_completed_
      -- 
    cp_elements(875) <= cp_elements(866);
    -- CP-element group 876 transition  bypass 
    -- predecessors 866 
    -- successors 873 
    -- members (4) 
      -- 	branch_block_stmt_2042/assign_stmt_3360_to_assign_stmt_3370/R_shifted_divisorx_x0x_xlcssax_xix_xix_xi_3363_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_3360_to_assign_stmt_3370/R_shifted_divisorx_x0x_xlcssax_xix_xix_xi_3363_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3360_to_assign_stmt_3370/R_shifted_divisorx_x0x_xlcssax_xix_xix_xi_3363_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_3360_to_assign_stmt_3370/R_shifted_divisorx_x0x_xlcssax_xix_xix_xi_3363_update_completed_
      -- 
    cp_elements(876) <= cp_elements(866);
    -- CP-element group 877 transition  input  bypass 
    -- predecessors 873 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_3360_to_assign_stmt_3370/SUB_u32_u32_3364_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3360_to_assign_stmt_3370/SUB_u32_u32_3364_Sample/$exit
      -- 	branch_block_stmt_2042/assign_stmt_3360_to_assign_stmt_3370/SUB_u32_u32_3364_Sample/ra
      -- 
    ra_13898_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => SUB_u32_u32_3364_inst_ack_0, ack => cp_elements(877)); -- 
    -- CP-element group 878 transition  input  bypass 
    -- predecessors 874 
    -- successors 879 
    -- members (7) 
      -- 	branch_block_stmt_2042/assign_stmt_3360_to_assign_stmt_3370/SUB_u32_u32_3364_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3360_to_assign_stmt_3370/SUB_u32_u32_3364_Update/$exit
      -- 	branch_block_stmt_2042/assign_stmt_3360_to_assign_stmt_3370/SUB_u32_u32_3364_Update/ca
      -- 	branch_block_stmt_2042/assign_stmt_3360_to_assign_stmt_3370/R_iNsTr_190_3367_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_3360_to_assign_stmt_3370/R_iNsTr_190_3367_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3360_to_assign_stmt_3370/R_iNsTr_190_3367_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_3360_to_assign_stmt_3370/R_iNsTr_190_3367_update_completed_
      -- 
    ca_13903_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => SUB_u32_u32_3364_inst_ack_1, ack => cp_elements(878)); -- 
    -- CP-element group 879 join  transition  output  bypass 
    -- predecessors 878 881 
    -- successors 882 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_3360_to_assign_stmt_3370/ULT_u32_u1_3369_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_3360_to_assign_stmt_3370/ULT_u32_u1_3369_Sample/$entry
      -- 	branch_block_stmt_2042/assign_stmt_3360_to_assign_stmt_3370/ULT_u32_u1_3369_Sample/rr
      -- 
    cp_element_group_879: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 20) := "cp_element_group_879"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(878) & cp_elements(881);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(879), clk => clk, reset => reset); --
    end block;
    rr_13919_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(879), ack => ULT_u32_u1_3369_inst_req_0); -- 
    -- CP-element group 880 transition  output  bypass 
    -- predecessors 866 
    -- successors 883 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_3360_to_assign_stmt_3370/ULT_u32_u1_3369_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_3360_to_assign_stmt_3370/ULT_u32_u1_3369_Update/$entry
      -- 	branch_block_stmt_2042/assign_stmt_3360_to_assign_stmt_3370/ULT_u32_u1_3369_Update/cr
      -- 
    cp_elements(880) <= cp_elements(866);
    cr_13924_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(880), ack => ULT_u32_u1_3369_inst_req_1); -- 
    -- CP-element group 881 transition  bypass 
    -- predecessors 866 
    -- successors 879 
    -- members (4) 
      -- 	branch_block_stmt_2042/assign_stmt_3360_to_assign_stmt_3370/R_iNsTr_97_3368_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_3360_to_assign_stmt_3370/R_iNsTr_97_3368_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3360_to_assign_stmt_3370/R_iNsTr_97_3368_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_3360_to_assign_stmt_3370/R_iNsTr_97_3368_update_completed_
      -- 
    cp_elements(881) <= cp_elements(866);
    -- CP-element group 882 transition  input  bypass 
    -- predecessors 879 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_3360_to_assign_stmt_3370/ULT_u32_u1_3369_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3360_to_assign_stmt_3370/ULT_u32_u1_3369_Sample/$exit
      -- 	branch_block_stmt_2042/assign_stmt_3360_to_assign_stmt_3370/ULT_u32_u1_3369_Sample/ra
      -- 
    ra_13920_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ULT_u32_u1_3369_inst_ack_0, ack => cp_elements(882)); -- 
    -- CP-element group 883 transition  input  bypass 
    -- predecessors 880 
    -- successors 884 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_3360_to_assign_stmt_3370/ULT_u32_u1_3369_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3360_to_assign_stmt_3370/ULT_u32_u1_3369_Update/$exit
      -- 	branch_block_stmt_2042/assign_stmt_3360_to_assign_stmt_3370/ULT_u32_u1_3369_Update/ca
      -- 
    ca_13925_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ULT_u32_u1_3369_inst_ack_1, ack => cp_elements(883)); -- 
    -- CP-element group 884 join  transition  bypass 
    -- predecessors 872 883 
    -- successors 53 
    -- members (1) 
      -- 	branch_block_stmt_2042/assign_stmt_3360_to_assign_stmt_3370/$exit
      -- 
    cp_element_group_884: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 20) := "cp_element_group_884"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(872) & cp_elements(883);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(884), clk => clk, reset => reset); --
    end block;
    -- CP-element group 885 transition  place  dead  bypass 
    -- predecessors 53 
    -- successors 54 
    -- members (8) 
      -- 	branch_block_stmt_2042/merge_stmt_3377__entry__
      -- 	branch_block_stmt_2042/if_stmt_3371__exit__
      -- 	branch_block_stmt_2042/if_stmt_3371_dead_link/$entry
      -- 	branch_block_stmt_2042/if_stmt_3371_dead_link/$exit
      -- 	branch_block_stmt_2042/if_stmt_3371_dead_link/dead_transition
      -- 	branch_block_stmt_2042/merge_stmt_3377_dead_link/$entry
      -- 	branch_block_stmt_2042/merge_stmt_3377_dead_link/$exit
      -- 	branch_block_stmt_2042/merge_stmt_3377_dead_link/dead_transition
      -- 
    cp_elements(885) <= false;
    -- CP-element group 886 transition  output  bypass 
    -- predecessors 53 
    -- successors 887 
    -- members (3) 
      -- 	branch_block_stmt_2042/if_stmt_3371_eval_test/$entry
      -- 	branch_block_stmt_2042/if_stmt_3371_eval_test/$exit
      -- 	branch_block_stmt_2042/if_stmt_3371_eval_test/branch_req
      -- 
    cp_elements(886) <= cp_elements(53);
    branch_req_13933_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(886), ack => if_stmt_3371_branch_req_0); -- 
    -- CP-element group 887 branch  place  bypass 
    -- predecessors 886 
    -- successors 888 890 
    -- members (1) 
      -- 	branch_block_stmt_2042/R_iNsTr_191_3372_place
      -- 
    cp_elements(887) <= cp_elements(886);
    -- CP-element group 888 transition  bypass 
    -- predecessors 887 
    -- successors 889 
    -- members (1) 
      -- 	branch_block_stmt_2042/if_stmt_3371_if_link/$entry
      -- 
    cp_elements(888) <= cp_elements(887);
    -- CP-element group 889 fork  transition  place  input  bypass 
    -- predecessors 888 
    -- successors 2130 2132 
    -- members (8) 
      -- 	branch_block_stmt_2042/if_stmt_3371_if_link/$exit
      -- 	branch_block_stmt_2042/if_stmt_3371_if_link/if_choice_transition
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi_xx_xloopexitx_xix_xix_xix_xloopexit
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi_xx_xloopexitx_xix_xix_xix_xloopexit_PhiReq/$entry
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi_xx_xloopexitx_xix_xix_xix_xloopexit_PhiReq/phi_stmt_3378/$entry
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi_xx_xloopexitx_xix_xix_xix_xloopexit_PhiReq/phi_stmt_3378/phi_stmt_3378_sources/$entry
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi_xx_xloopexitx_xix_xix_xix_xloopexit_PhiReq/phi_stmt_3378/phi_stmt_3378_sources/type_cast_3381/$entry
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi_xx_xloopexitx_xix_xix_xix_xloopexit_PhiReq/phi_stmt_3378/phi_stmt_3378_sources/type_cast_3381/SplitProtocol/$entry
      -- 
    if_choice_transition_13938_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_3371_branch_ack_1, ack => cp_elements(889)); -- 
    -- CP-element group 890 transition  bypass 
    -- predecessors 887 
    -- successors 891 
    -- members (1) 
      -- 	branch_block_stmt_2042/if_stmt_3371_else_link/$entry
      -- 
    cp_elements(890) <= cp_elements(887);
    -- CP-element group 891 transition  place  input  bypass 
    -- predecessors 890 
    -- successors 2000 
    -- members (3) 
      -- 	branch_block_stmt_2042/if_stmt_3371_else_link/$exit
      -- 	branch_block_stmt_2042/if_stmt_3371_else_link/else_choice_transition
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi_bbx_xnph7x_xix_xix_xi
      -- 
    else_choice_transition_13942_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_3371_branch_ack_0, ack => cp_elements(891)); -- 
    -- CP-element group 892 fork  transition  bypass 
    -- predecessors 2171 
    -- successors 893 894 897 900 901 907 
    -- members (1) 
      -- 	branch_block_stmt_2042/assign_stmt_3407_to_assign_stmt_3426/$entry
      -- 
    cp_elements(892) <= cp_elements(2171);
    -- CP-element group 893 transition  output  bypass 
    -- predecessors 892 
    -- successors 896 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_3407_to_assign_stmt_3426/AND_u32_u32_3406_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_3407_to_assign_stmt_3426/AND_u32_u32_3406_Update/$entry
      -- 	branch_block_stmt_2042/assign_stmt_3407_to_assign_stmt_3426/AND_u32_u32_3406_Update/cr
      -- 
    cp_elements(893) <= cp_elements(892);
    cr_13964_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(893), ack => AND_u32_u32_3406_inst_req_1); -- 
    -- CP-element group 894 transition  output  bypass 
    -- predecessors 892 
    -- successors 895 
    -- members (7) 
      -- 	branch_block_stmt_2042/assign_stmt_3407_to_assign_stmt_3426/AND_u32_u32_3406_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_3407_to_assign_stmt_3426/R_tempx_x0x_xphx_xix_xi_3403_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_3407_to_assign_stmt_3426/R_tempx_x0x_xphx_xix_xi_3403_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3407_to_assign_stmt_3426/R_tempx_x0x_xphx_xix_xi_3403_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_3407_to_assign_stmt_3426/R_tempx_x0x_xphx_xix_xi_3403_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3407_to_assign_stmt_3426/AND_u32_u32_3406_Sample/$entry
      -- 	branch_block_stmt_2042/assign_stmt_3407_to_assign_stmt_3426/AND_u32_u32_3406_Sample/rr
      -- 
    cp_elements(894) <= cp_elements(892);
    rr_13959_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(894), ack => AND_u32_u32_3406_inst_req_0); -- 
    -- CP-element group 895 transition  input  bypass 
    -- predecessors 894 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_3407_to_assign_stmt_3426/AND_u32_u32_3406_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3407_to_assign_stmt_3426/AND_u32_u32_3406_Sample/$exit
      -- 	branch_block_stmt_2042/assign_stmt_3407_to_assign_stmt_3426/AND_u32_u32_3406_Sample/ra
      -- 
    ra_13960_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => AND_u32_u32_3406_inst_ack_0, ack => cp_elements(895)); -- 
    -- CP-element group 896 transition  input  output  bypass 
    -- predecessors 893 
    -- successors 898 
    -- members (10) 
      -- 	branch_block_stmt_2042/assign_stmt_3407_to_assign_stmt_3426/AND_u32_u32_3406_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3407_to_assign_stmt_3426/AND_u32_u32_3406_Update/$exit
      -- 	branch_block_stmt_2042/assign_stmt_3407_to_assign_stmt_3426/AND_u32_u32_3406_Update/ca
      -- 	branch_block_stmt_2042/assign_stmt_3407_to_assign_stmt_3426/EQ_u32_u1_3412_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_3407_to_assign_stmt_3426/R_iNsTr_121_3409_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_3407_to_assign_stmt_3426/R_iNsTr_121_3409_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3407_to_assign_stmt_3426/R_iNsTr_121_3409_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_3407_to_assign_stmt_3426/R_iNsTr_121_3409_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3407_to_assign_stmt_3426/EQ_u32_u1_3412_Sample/$entry
      -- 	branch_block_stmt_2042/assign_stmt_3407_to_assign_stmt_3426/EQ_u32_u1_3412_Sample/rr
      -- 
    ca_13965_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => AND_u32_u32_3406_inst_ack_1, ack => cp_elements(896)); -- 
    rr_13977_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(896), ack => EQ_u32_u1_3412_inst_req_0); -- 
    -- CP-element group 897 transition  output  bypass 
    -- predecessors 892 
    -- successors 899 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_3407_to_assign_stmt_3426/EQ_u32_u1_3412_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_3407_to_assign_stmt_3426/EQ_u32_u1_3412_Update/$entry
      -- 	branch_block_stmt_2042/assign_stmt_3407_to_assign_stmt_3426/EQ_u32_u1_3412_Update/cr
      -- 
    cp_elements(897) <= cp_elements(892);
    cr_13982_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(897), ack => EQ_u32_u1_3412_inst_req_1); -- 
    -- CP-element group 898 transition  input  bypass 
    -- predecessors 896 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_3407_to_assign_stmt_3426/EQ_u32_u1_3412_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3407_to_assign_stmt_3426/EQ_u32_u1_3412_Sample/$exit
      -- 	branch_block_stmt_2042/assign_stmt_3407_to_assign_stmt_3426/EQ_u32_u1_3412_Sample/ra
      -- 
    ra_13978_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u32_u1_3412_inst_ack_0, ack => cp_elements(898)); -- 
    -- CP-element group 899 transition  input  bypass 
    -- predecessors 897 
    -- successors 906 
    -- members (7) 
      -- 	branch_block_stmt_2042/assign_stmt_3407_to_assign_stmt_3426/EQ_u32_u1_3412_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3407_to_assign_stmt_3426/EQ_u32_u1_3412_Update/$exit
      -- 	branch_block_stmt_2042/assign_stmt_3407_to_assign_stmt_3426/EQ_u32_u1_3412_Update/ca
      -- 	branch_block_stmt_2042/assign_stmt_3407_to_assign_stmt_3426/R_iNsTr_122_3423_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_3407_to_assign_stmt_3426/R_iNsTr_122_3423_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3407_to_assign_stmt_3426/R_iNsTr_122_3423_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_3407_to_assign_stmt_3426/R_iNsTr_122_3423_update_completed_
      -- 
    ca_13983_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u32_u1_3412_inst_ack_1, ack => cp_elements(899)); -- 
    -- CP-element group 900 transition  output  bypass 
    -- predecessors 892 
    -- successors 905 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_3407_to_assign_stmt_3426/NEQ_i32_u1_3420_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_3407_to_assign_stmt_3426/NEQ_i32_u1_3420_Update/$entry
      -- 	branch_block_stmt_2042/assign_stmt_3407_to_assign_stmt_3426/NEQ_i32_u1_3420_Update/cr
      -- 
    cp_elements(900) <= cp_elements(892);
    cr_14014_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(900), ack => NEQ_i32_u1_3420_inst_req_1); -- 
    -- CP-element group 901 transition  output  bypass 
    -- predecessors 892 
    -- successors 902 
    -- members (7) 
      -- 	branch_block_stmt_2042/assign_stmt_3407_to_assign_stmt_3426/type_cast_3416_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_3407_to_assign_stmt_3426/R_tempx_x0x_xphx_xix_xi_3415_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_3407_to_assign_stmt_3426/R_tempx_x0x_xphx_xix_xi_3415_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3407_to_assign_stmt_3426/R_tempx_x0x_xphx_xix_xi_3415_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_3407_to_assign_stmt_3426/R_tempx_x0x_xphx_xix_xi_3415_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3407_to_assign_stmt_3426/type_cast_3416_Sample/$entry
      -- 	branch_block_stmt_2042/assign_stmt_3407_to_assign_stmt_3426/type_cast_3416_Sample/rr
      -- 
    cp_elements(901) <= cp_elements(892);
    rr_13999_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(901), ack => type_cast_3416_inst_req_0); -- 
    -- CP-element group 902 transition  input  output  bypass 
    -- predecessors 901 
    -- successors 903 
    -- members (6) 
      -- 	branch_block_stmt_2042/assign_stmt_3407_to_assign_stmt_3426/type_cast_3416_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3407_to_assign_stmt_3426/type_cast_3416_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_3407_to_assign_stmt_3426/type_cast_3416_Sample/$exit
      -- 	branch_block_stmt_2042/assign_stmt_3407_to_assign_stmt_3426/type_cast_3416_Sample/ra
      -- 	branch_block_stmt_2042/assign_stmt_3407_to_assign_stmt_3426/type_cast_3416_Update/$entry
      -- 	branch_block_stmt_2042/assign_stmt_3407_to_assign_stmt_3426/type_cast_3416_Update/cr
      -- 
    ra_14000_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3416_inst_ack_0, ack => cp_elements(902)); -- 
    cr_14004_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(902), ack => type_cast_3416_inst_req_1); -- 
    -- CP-element group 903 transition  input  output  bypass 
    -- predecessors 902 
    -- successors 904 
    -- members (6) 
      -- 	branch_block_stmt_2042/assign_stmt_3407_to_assign_stmt_3426/NEQ_i32_u1_3420_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_3407_to_assign_stmt_3426/type_cast_3416_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3407_to_assign_stmt_3426/type_cast_3416_Update/$exit
      -- 	branch_block_stmt_2042/assign_stmt_3407_to_assign_stmt_3426/type_cast_3416_Update/ca
      -- 	branch_block_stmt_2042/assign_stmt_3407_to_assign_stmt_3426/NEQ_i32_u1_3420_Sample/$entry
      -- 	branch_block_stmt_2042/assign_stmt_3407_to_assign_stmt_3426/NEQ_i32_u1_3420_Sample/rr
      -- 
    ca_14005_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3416_inst_ack_1, ack => cp_elements(903)); -- 
    rr_14009_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(903), ack => NEQ_i32_u1_3420_inst_req_0); -- 
    -- CP-element group 904 transition  input  bypass 
    -- predecessors 903 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_3407_to_assign_stmt_3426/NEQ_i32_u1_3420_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3407_to_assign_stmt_3426/NEQ_i32_u1_3420_Sample/$exit
      -- 	branch_block_stmt_2042/assign_stmt_3407_to_assign_stmt_3426/NEQ_i32_u1_3420_Sample/ra
      -- 
    ra_14010_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => NEQ_i32_u1_3420_inst_ack_0, ack => cp_elements(904)); -- 
    -- CP-element group 905 transition  input  bypass 
    -- predecessors 900 
    -- successors 906 
    -- members (7) 
      -- 	branch_block_stmt_2042/assign_stmt_3407_to_assign_stmt_3426/NEQ_i32_u1_3420_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3407_to_assign_stmt_3426/NEQ_i32_u1_3420_Update/$exit
      -- 	branch_block_stmt_2042/assign_stmt_3407_to_assign_stmt_3426/NEQ_i32_u1_3420_Update/ca
      -- 	branch_block_stmt_2042/assign_stmt_3407_to_assign_stmt_3426/R_iNsTr_123_3424_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_3407_to_assign_stmt_3426/R_iNsTr_123_3424_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3407_to_assign_stmt_3426/R_iNsTr_123_3424_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_3407_to_assign_stmt_3426/R_iNsTr_123_3424_update_completed_
      -- 
    ca_14015_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => NEQ_i32_u1_3420_inst_ack_1, ack => cp_elements(905)); -- 
    -- CP-element group 906 join  transition  output  bypass 
    -- predecessors 899 905 
    -- successors 908 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_3407_to_assign_stmt_3426/AND_u1_u1_3425_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_3407_to_assign_stmt_3426/AND_u1_u1_3425_Sample/$entry
      -- 	branch_block_stmt_2042/assign_stmt_3407_to_assign_stmt_3426/AND_u1_u1_3425_Sample/rr
      -- 
    cp_element_group_906: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 20) := "cp_element_group_906"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(899) & cp_elements(905);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(906), clk => clk, reset => reset); --
    end block;
    rr_14031_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(906), ack => AND_u1_u1_3425_inst_req_0); -- 
    -- CP-element group 907 transition  output  bypass 
    -- predecessors 892 
    -- successors 909 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_3407_to_assign_stmt_3426/AND_u1_u1_3425_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_3407_to_assign_stmt_3426/AND_u1_u1_3425_Update/$entry
      -- 	branch_block_stmt_2042/assign_stmt_3407_to_assign_stmt_3426/AND_u1_u1_3425_Update/cr
      -- 
    cp_elements(907) <= cp_elements(892);
    cr_14036_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(907), ack => AND_u1_u1_3425_inst_req_1); -- 
    -- CP-element group 908 transition  input  bypass 
    -- predecessors 906 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_3407_to_assign_stmt_3426/AND_u1_u1_3425_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3407_to_assign_stmt_3426/AND_u1_u1_3425_Sample/$exit
      -- 	branch_block_stmt_2042/assign_stmt_3407_to_assign_stmt_3426/AND_u1_u1_3425_Sample/ra
      -- 
    ra_14032_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => AND_u1_u1_3425_inst_ack_0, ack => cp_elements(908)); -- 
    -- CP-element group 909 branch  transition  place  input  bypass 
    -- predecessors 907 
    -- successors 910 911 
    -- members (6) 
      -- 	branch_block_stmt_2042/if_stmt_3427__entry__
      -- 	branch_block_stmt_2042/assign_stmt_3407_to_assign_stmt_3426__exit__
      -- 	branch_block_stmt_2042/assign_stmt_3407_to_assign_stmt_3426/$exit
      -- 	branch_block_stmt_2042/assign_stmt_3407_to_assign_stmt_3426/AND_u1_u1_3425_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3407_to_assign_stmt_3426/AND_u1_u1_3425_Update/$exit
      -- 	branch_block_stmt_2042/assign_stmt_3407_to_assign_stmt_3426/AND_u1_u1_3425_Update/ca
      -- 
    ca_14037_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => AND_u1_u1_3425_inst_ack_1, ack => cp_elements(909)); -- 
    -- CP-element group 910 transition  place  dead  bypass 
    -- predecessors 909 
    -- successors 55 
    -- members (8) 
      -- 	branch_block_stmt_2042/merge_stmt_3433__entry__
      -- 	branch_block_stmt_2042/if_stmt_3427__exit__
      -- 	branch_block_stmt_2042/if_stmt_3427_dead_link/$entry
      -- 	branch_block_stmt_2042/if_stmt_3427_dead_link/$exit
      -- 	branch_block_stmt_2042/if_stmt_3427_dead_link/dead_transition
      -- 	branch_block_stmt_2042/merge_stmt_3433_dead_link/dead_transition
      -- 	branch_block_stmt_2042/merge_stmt_3433_dead_link/$exit
      -- 	branch_block_stmt_2042/merge_stmt_3433_dead_link/$entry
      -- 
    cp_elements(910) <= false;
    -- CP-element group 911 transition  output  bypass 
    -- predecessors 909 
    -- successors 912 
    -- members (3) 
      -- 	branch_block_stmt_2042/if_stmt_3427_eval_test/$entry
      -- 	branch_block_stmt_2042/if_stmt_3427_eval_test/$exit
      -- 	branch_block_stmt_2042/if_stmt_3427_eval_test/branch_req
      -- 
    cp_elements(911) <= cp_elements(909);
    branch_req_14045_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(911), ack => if_stmt_3427_branch_req_0); -- 
    -- CP-element group 912 branch  place  bypass 
    -- predecessors 911 
    -- successors 913 915 
    -- members (1) 
      -- 	branch_block_stmt_2042/R_orx_xcond11x_xix_xi_3428_place
      -- 
    cp_elements(912) <= cp_elements(911);
    -- CP-element group 913 transition  bypass 
    -- predecessors 912 
    -- successors 914 
    -- members (1) 
      -- 	branch_block_stmt_2042/if_stmt_3427_if_link/$entry
      -- 
    cp_elements(913) <= cp_elements(912);
    -- CP-element group 914 transition  place  input  bypass 
    -- predecessors 913 
    -- successors 55 
    -- members (9) 
      -- 	branch_block_stmt_2042/if_stmt_3427_if_link/$exit
      -- 	branch_block_stmt_2042/if_stmt_3427_if_link/if_choice_transition
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xpreheaderx_xix_xi_udiv32x_xexitx_xix_xix_xpreheader
      -- 	branch_block_stmt_2042/merge_stmt_3433_PhiAck/dummy
      -- 	branch_block_stmt_2042/merge_stmt_3433_PhiAck/$exit
      -- 	branch_block_stmt_2042/merge_stmt_3433_PhiAck/$entry
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xpreheaderx_xix_xi_udiv32x_xexitx_xix_xix_xpreheader_PhiReq/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xpreheaderx_xix_xi_udiv32x_xexitx_xix_xix_xpreheader_PhiReq/$entry
      -- 	branch_block_stmt_2042/merge_stmt_3433_PhiReqMerge
      -- 
    if_choice_transition_14050_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_3427_branch_ack_1, ack => cp_elements(914)); -- 
    -- CP-element group 915 transition  bypass 
    -- predecessors 912 
    -- successors 916 
    -- members (1) 
      -- 	branch_block_stmt_2042/if_stmt_3427_else_link/$entry
      -- 
    cp_elements(915) <= cp_elements(912);
    -- CP-element group 916 transition  place  input  bypass 
    -- predecessors 915 
    -- successors 2234 
    -- members (3) 
      -- 	branch_block_stmt_2042/if_stmt_3427_else_link/$exit
      -- 	branch_block_stmt_2042/if_stmt_3427_else_link/else_choice_transition
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xpreheaderx_xix_xi_xx_xcritedgex_xix_xi
      -- 
    else_choice_transition_14054_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_3427_branch_ack_0, ack => cp_elements(916)); -- 
    -- CP-element group 917 fork  transition  bypass 
    -- predecessors 56 
    -- successors 918 919 922 926 929 936 939 940 
    -- members (1) 
      -- 	branch_block_stmt_2042/assign_stmt_3455_to_assign_stmt_3486/$entry
      -- 
    cp_elements(917) <= cp_elements(56);
    -- CP-element group 918 transition  output  bypass 
    -- predecessors 917 
    -- successors 921 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_3455_to_assign_stmt_3486/SHL_u32_u32_3454_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_3455_to_assign_stmt_3486/SHL_u32_u32_3454_Update/$entry
      -- 	branch_block_stmt_2042/assign_stmt_3455_to_assign_stmt_3486/SHL_u32_u32_3454_Update/cr
      -- 
    cp_elements(918) <= cp_elements(917);
    cr_14076_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(918), ack => SHL_u32_u32_3454_inst_req_1); -- 
    -- CP-element group 919 transition  output  bypass 
    -- predecessors 917 
    -- successors 920 
    -- members (7) 
      -- 	branch_block_stmt_2042/assign_stmt_3455_to_assign_stmt_3486/SHL_u32_u32_3454_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_3455_to_assign_stmt_3486/R_tempx_x012x_xix_xi_3451_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_3455_to_assign_stmt_3486/R_tempx_x012x_xix_xi_3451_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3455_to_assign_stmt_3486/R_tempx_x012x_xix_xi_3451_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_3455_to_assign_stmt_3486/R_tempx_x012x_xix_xi_3451_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3455_to_assign_stmt_3486/SHL_u32_u32_3454_Sample/$entry
      -- 	branch_block_stmt_2042/assign_stmt_3455_to_assign_stmt_3486/SHL_u32_u32_3454_Sample/rr
      -- 
    cp_elements(919) <= cp_elements(917);
    rr_14071_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(919), ack => SHL_u32_u32_3454_inst_req_0); -- 
    -- CP-element group 920 transition  input  bypass 
    -- predecessors 919 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_3455_to_assign_stmt_3486/SHL_u32_u32_3454_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3455_to_assign_stmt_3486/SHL_u32_u32_3454_Sample/$exit
      -- 	branch_block_stmt_2042/assign_stmt_3455_to_assign_stmt_3486/SHL_u32_u32_3454_Sample/ra
      -- 
    ra_14072_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => SHL_u32_u32_3454_inst_ack_0, ack => cp_elements(920)); -- 
    -- CP-element group 921 fork  transition  input  bypass 
    -- predecessors 918 
    -- successors 923 930 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_3455_to_assign_stmt_3486/SHL_u32_u32_3454_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3455_to_assign_stmt_3486/SHL_u32_u32_3454_Update/$exit
      -- 	branch_block_stmt_2042/assign_stmt_3455_to_assign_stmt_3486/SHL_u32_u32_3454_Update/ca
      -- 
    ca_14077_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => SHL_u32_u32_3454_inst_ack_1, ack => cp_elements(921)); -- 
    -- CP-element group 922 transition  output  bypass 
    -- predecessors 917 
    -- successors 925 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_3455_to_assign_stmt_3486/AND_u32_u32_3460_Update/cr
      -- 	branch_block_stmt_2042/assign_stmt_3455_to_assign_stmt_3486/AND_u32_u32_3460_Update/$entry
      -- 	branch_block_stmt_2042/assign_stmt_3455_to_assign_stmt_3486/AND_u32_u32_3460_update_start_
      -- 
    cp_elements(922) <= cp_elements(917);
    cr_14094_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(922), ack => AND_u32_u32_3460_inst_req_1); -- 
    -- CP-element group 923 transition  output  bypass 
    -- predecessors 921 
    -- successors 924 
    -- members (7) 
      -- 	branch_block_stmt_2042/assign_stmt_3455_to_assign_stmt_3486/AND_u32_u32_3460_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_3455_to_assign_stmt_3486/R_iNsTr_194_3457_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_3455_to_assign_stmt_3486/R_iNsTr_194_3457_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3455_to_assign_stmt_3486/R_iNsTr_194_3457_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_3455_to_assign_stmt_3486/R_iNsTr_194_3457_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3455_to_assign_stmt_3486/AND_u32_u32_3460_Sample/$entry
      -- 	branch_block_stmt_2042/assign_stmt_3455_to_assign_stmt_3486/AND_u32_u32_3460_Sample/rr
      -- 
    cp_elements(923) <= cp_elements(921);
    rr_14089_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(923), ack => AND_u32_u32_3460_inst_req_0); -- 
    -- CP-element group 924 transition  input  bypass 
    -- predecessors 923 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_3455_to_assign_stmt_3486/AND_u32_u32_3460_Sample/ra
      -- 	branch_block_stmt_2042/assign_stmt_3455_to_assign_stmt_3486/AND_u32_u32_3460_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3455_to_assign_stmt_3486/AND_u32_u32_3460_Sample/$exit
      -- 
    ra_14090_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => AND_u32_u32_3460_inst_ack_0, ack => cp_elements(924)); -- 
    -- CP-element group 925 transition  input  output  bypass 
    -- predecessors 922 
    -- successors 927 
    -- members (10) 
      -- 	branch_block_stmt_2042/assign_stmt_3455_to_assign_stmt_3486/AND_u32_u32_3460_Update/ca
      -- 	branch_block_stmt_2042/assign_stmt_3455_to_assign_stmt_3486/EQ_u32_u1_3466_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_3455_to_assign_stmt_3486/R_iNsTr_195_3463_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3455_to_assign_stmt_3486/AND_u32_u32_3460_Update/$exit
      -- 	branch_block_stmt_2042/assign_stmt_3455_to_assign_stmt_3486/R_iNsTr_195_3463_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_3455_to_assign_stmt_3486/R_iNsTr_195_3463_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_3455_to_assign_stmt_3486/R_iNsTr_195_3463_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3455_to_assign_stmt_3486/AND_u32_u32_3460_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3455_to_assign_stmt_3486/EQ_u32_u1_3466_Sample/$entry
      -- 	branch_block_stmt_2042/assign_stmt_3455_to_assign_stmt_3486/EQ_u32_u1_3466_Sample/rr
      -- 
    ca_14095_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => AND_u32_u32_3460_inst_ack_1, ack => cp_elements(925)); -- 
    rr_14107_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(925), ack => EQ_u32_u1_3466_inst_req_0); -- 
    -- CP-element group 926 transition  output  bypass 
    -- predecessors 917 
    -- successors 928 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_3455_to_assign_stmt_3486/EQ_u32_u1_3466_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_3455_to_assign_stmt_3486/EQ_u32_u1_3466_Update/$entry
      -- 	branch_block_stmt_2042/assign_stmt_3455_to_assign_stmt_3486/EQ_u32_u1_3466_Update/cr
      -- 
    cp_elements(926) <= cp_elements(917);
    cr_14112_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(926), ack => EQ_u32_u1_3466_inst_req_1); -- 
    -- CP-element group 927 transition  input  bypass 
    -- predecessors 925 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_3455_to_assign_stmt_3486/EQ_u32_u1_3466_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3455_to_assign_stmt_3486/EQ_u32_u1_3466_Sample/$exit
      -- 	branch_block_stmt_2042/assign_stmt_3455_to_assign_stmt_3486/EQ_u32_u1_3466_Sample/ra
      -- 
    ra_14108_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u32_u1_3466_inst_ack_0, ack => cp_elements(927)); -- 
    -- CP-element group 928 transition  input  bypass 
    -- predecessors 926 
    -- successors 935 
    -- members (7) 
      -- 	branch_block_stmt_2042/assign_stmt_3455_to_assign_stmt_3486/EQ_u32_u1_3466_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3455_to_assign_stmt_3486/EQ_u32_u1_3466_Update/$exit
      -- 	branch_block_stmt_2042/assign_stmt_3455_to_assign_stmt_3486/EQ_u32_u1_3466_Update/ca
      -- 	branch_block_stmt_2042/assign_stmt_3455_to_assign_stmt_3486/R_iNsTr_196_3477_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_3455_to_assign_stmt_3486/R_iNsTr_196_3477_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3455_to_assign_stmt_3486/R_iNsTr_196_3477_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_3455_to_assign_stmt_3486/R_iNsTr_196_3477_update_completed_
      -- 
    ca_14113_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u32_u1_3466_inst_ack_1, ack => cp_elements(928)); -- 
    -- CP-element group 929 transition  output  bypass 
    -- predecessors 917 
    -- successors 934 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_3455_to_assign_stmt_3486/NEQ_i32_u1_3474_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_3455_to_assign_stmt_3486/NEQ_i32_u1_3474_Update/$entry
      -- 	branch_block_stmt_2042/assign_stmt_3455_to_assign_stmt_3486/NEQ_i32_u1_3474_Update/cr
      -- 
    cp_elements(929) <= cp_elements(917);
    cr_14144_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(929), ack => NEQ_i32_u1_3474_inst_req_1); -- 
    -- CP-element group 930 transition  output  bypass 
    -- predecessors 921 
    -- successors 931 
    -- members (7) 
      -- 	branch_block_stmt_2042/assign_stmt_3455_to_assign_stmt_3486/type_cast_3470_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_3455_to_assign_stmt_3486/R_iNsTr_194_3469_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_3455_to_assign_stmt_3486/R_iNsTr_194_3469_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3455_to_assign_stmt_3486/R_iNsTr_194_3469_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_3455_to_assign_stmt_3486/R_iNsTr_194_3469_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3455_to_assign_stmt_3486/type_cast_3470_Sample/$entry
      -- 	branch_block_stmt_2042/assign_stmt_3455_to_assign_stmt_3486/type_cast_3470_Sample/rr
      -- 
    cp_elements(930) <= cp_elements(921);
    rr_14129_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(930), ack => type_cast_3470_inst_req_0); -- 
    -- CP-element group 931 transition  input  output  bypass 
    -- predecessors 930 
    -- successors 932 
    -- members (6) 
      -- 	branch_block_stmt_2042/assign_stmt_3455_to_assign_stmt_3486/type_cast_3470_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3455_to_assign_stmt_3486/type_cast_3470_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_3455_to_assign_stmt_3486/type_cast_3470_Sample/$exit
      -- 	branch_block_stmt_2042/assign_stmt_3455_to_assign_stmt_3486/type_cast_3470_Sample/ra
      -- 	branch_block_stmt_2042/assign_stmt_3455_to_assign_stmt_3486/type_cast_3470_Update/$entry
      -- 	branch_block_stmt_2042/assign_stmt_3455_to_assign_stmt_3486/type_cast_3470_Update/cr
      -- 
    ra_14130_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3470_inst_ack_0, ack => cp_elements(931)); -- 
    cr_14134_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(931), ack => type_cast_3470_inst_req_1); -- 
    -- CP-element group 932 transition  input  output  bypass 
    -- predecessors 931 
    -- successors 933 
    -- members (6) 
      -- 	branch_block_stmt_2042/assign_stmt_3455_to_assign_stmt_3486/NEQ_i32_u1_3474_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_3455_to_assign_stmt_3486/type_cast_3470_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3455_to_assign_stmt_3486/type_cast_3470_Update/$exit
      -- 	branch_block_stmt_2042/assign_stmt_3455_to_assign_stmt_3486/type_cast_3470_Update/ca
      -- 	branch_block_stmt_2042/assign_stmt_3455_to_assign_stmt_3486/NEQ_i32_u1_3474_Sample/$entry
      -- 	branch_block_stmt_2042/assign_stmt_3455_to_assign_stmt_3486/NEQ_i32_u1_3474_Sample/rr
      -- 
    ca_14135_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3470_inst_ack_1, ack => cp_elements(932)); -- 
    rr_14139_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(932), ack => NEQ_i32_u1_3474_inst_req_0); -- 
    -- CP-element group 933 transition  input  bypass 
    -- predecessors 932 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_3455_to_assign_stmt_3486/NEQ_i32_u1_3474_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3455_to_assign_stmt_3486/NEQ_i32_u1_3474_Sample/$exit
      -- 	branch_block_stmt_2042/assign_stmt_3455_to_assign_stmt_3486/NEQ_i32_u1_3474_Sample/ra
      -- 
    ra_14140_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => NEQ_i32_u1_3474_inst_ack_0, ack => cp_elements(933)); -- 
    -- CP-element group 934 transition  input  bypass 
    -- predecessors 929 
    -- successors 935 
    -- members (7) 
      -- 	branch_block_stmt_2042/assign_stmt_3455_to_assign_stmt_3486/NEQ_i32_u1_3474_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3455_to_assign_stmt_3486/NEQ_i32_u1_3474_Update/$exit
      -- 	branch_block_stmt_2042/assign_stmt_3455_to_assign_stmt_3486/NEQ_i32_u1_3474_Update/ca
      -- 	branch_block_stmt_2042/assign_stmt_3455_to_assign_stmt_3486/R_iNsTr_197_3478_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_3455_to_assign_stmt_3486/R_iNsTr_197_3478_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3455_to_assign_stmt_3486/R_iNsTr_197_3478_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_3455_to_assign_stmt_3486/R_iNsTr_197_3478_update_completed_
      -- 
    ca_14145_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => NEQ_i32_u1_3474_inst_ack_1, ack => cp_elements(934)); -- 
    -- CP-element group 935 join  transition  output  bypass 
    -- predecessors 928 934 
    -- successors 937 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_3455_to_assign_stmt_3486/AND_u1_u1_3479_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_3455_to_assign_stmt_3486/AND_u1_u1_3479_Sample/$entry
      -- 	branch_block_stmt_2042/assign_stmt_3455_to_assign_stmt_3486/AND_u1_u1_3479_Sample/rr
      -- 
    cp_element_group_935: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 20) := "cp_element_group_935"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(928) & cp_elements(934);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(935), clk => clk, reset => reset); --
    end block;
    rr_14161_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(935), ack => AND_u1_u1_3479_inst_req_0); -- 
    -- CP-element group 936 transition  output  bypass 
    -- predecessors 917 
    -- successors 938 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_3455_to_assign_stmt_3486/AND_u1_u1_3479_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_3455_to_assign_stmt_3486/AND_u1_u1_3479_Update/$entry
      -- 	branch_block_stmt_2042/assign_stmt_3455_to_assign_stmt_3486/AND_u1_u1_3479_Update/cr
      -- 
    cp_elements(936) <= cp_elements(917);
    cr_14166_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(936), ack => AND_u1_u1_3479_inst_req_1); -- 
    -- CP-element group 937 transition  input  bypass 
    -- predecessors 935 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_3455_to_assign_stmt_3486/AND_u1_u1_3479_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3455_to_assign_stmt_3486/AND_u1_u1_3479_Sample/$exit
      -- 	branch_block_stmt_2042/assign_stmt_3455_to_assign_stmt_3486/AND_u1_u1_3479_Sample/ra
      -- 
    ra_14162_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => AND_u1_u1_3479_inst_ack_0, ack => cp_elements(937)); -- 
    -- CP-element group 938 transition  input  bypass 
    -- predecessors 936 
    -- successors 943 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_3455_to_assign_stmt_3486/AND_u1_u1_3479_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3455_to_assign_stmt_3486/AND_u1_u1_3479_Update/$exit
      -- 	branch_block_stmt_2042/assign_stmt_3455_to_assign_stmt_3486/AND_u1_u1_3479_Update/ca
      -- 
    ca_14167_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => AND_u1_u1_3479_inst_ack_1, ack => cp_elements(938)); -- 
    -- CP-element group 939 transition  output  bypass 
    -- predecessors 917 
    -- successors 942 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_3455_to_assign_stmt_3486/ADD_u32_u32_3485_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_3455_to_assign_stmt_3486/ADD_u32_u32_3485_Update/$entry
      -- 	branch_block_stmt_2042/assign_stmt_3455_to_assign_stmt_3486/ADD_u32_u32_3485_Update/cr
      -- 
    cp_elements(939) <= cp_elements(917);
    cr_14184_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(939), ack => ADD_u32_u32_3485_inst_req_1); -- 
    -- CP-element group 940 transition  output  bypass 
    -- predecessors 917 
    -- successors 941 
    -- members (7) 
      -- 	branch_block_stmt_2042/assign_stmt_3455_to_assign_stmt_3486/R_iNsTr_193_3482_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3455_to_assign_stmt_3486/ADD_u32_u32_3485_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_3455_to_assign_stmt_3486/R_iNsTr_193_3482_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_3455_to_assign_stmt_3486/R_iNsTr_193_3482_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_3455_to_assign_stmt_3486/R_iNsTr_193_3482_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3455_to_assign_stmt_3486/ADD_u32_u32_3485_Sample/$entry
      -- 	branch_block_stmt_2042/assign_stmt_3455_to_assign_stmt_3486/ADD_u32_u32_3485_Sample/rr
      -- 
    cp_elements(940) <= cp_elements(917);
    rr_14179_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(940), ack => ADD_u32_u32_3485_inst_req_0); -- 
    -- CP-element group 941 transition  input  bypass 
    -- predecessors 940 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_3455_to_assign_stmt_3486/ADD_u32_u32_3485_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3455_to_assign_stmt_3486/ADD_u32_u32_3485_Sample/$exit
      -- 	branch_block_stmt_2042/assign_stmt_3455_to_assign_stmt_3486/ADD_u32_u32_3485_Sample/ra
      -- 
    ra_14180_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u32_u32_3485_inst_ack_0, ack => cp_elements(941)); -- 
    -- CP-element group 942 transition  input  bypass 
    -- predecessors 939 
    -- successors 943 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_3455_to_assign_stmt_3486/ADD_u32_u32_3485_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3455_to_assign_stmt_3486/ADD_u32_u32_3485_Update/$exit
      -- 	branch_block_stmt_2042/assign_stmt_3455_to_assign_stmt_3486/ADD_u32_u32_3485_Update/ca
      -- 
    ca_14185_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u32_u32_3485_inst_ack_1, ack => cp_elements(942)); -- 
    -- CP-element group 943 join  transition  bypass 
    -- predecessors 938 942 
    -- successors 57 
    -- members (1) 
      -- 	branch_block_stmt_2042/assign_stmt_3455_to_assign_stmt_3486/$exit
      -- 
    cp_element_group_943: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 20) := "cp_element_group_943"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(938) & cp_elements(942);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(943), clk => clk, reset => reset); --
    end block;
    -- CP-element group 944 transition  place  dead  bypass 
    -- predecessors 57 
    -- successors 58 
    -- members (8) 
      -- 	branch_block_stmt_2042/merge_stmt_3493__entry__
      -- 	branch_block_stmt_2042/if_stmt_3487__exit__
      -- 	branch_block_stmt_2042/if_stmt_3487_dead_link/$entry
      -- 	branch_block_stmt_2042/if_stmt_3487_dead_link/$exit
      -- 	branch_block_stmt_2042/if_stmt_3487_dead_link/dead_transition
      -- 	branch_block_stmt_2042/merge_stmt_3493_dead_link/$entry
      -- 	branch_block_stmt_2042/merge_stmt_3493_dead_link/$exit
      -- 	branch_block_stmt_2042/merge_stmt_3493_dead_link/dead_transition
      -- 
    cp_elements(944) <= false;
    -- CP-element group 945 transition  output  bypass 
    -- predecessors 57 
    -- successors 946 
    -- members (3) 
      -- 	branch_block_stmt_2042/if_stmt_3487_eval_test/$entry
      -- 	branch_block_stmt_2042/if_stmt_3487_eval_test/$exit
      -- 	branch_block_stmt_2042/if_stmt_3487_eval_test/branch_req
      -- 
    cp_elements(945) <= cp_elements(57);
    branch_req_14193_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(945), ack => if_stmt_3487_branch_req_0); -- 
    -- CP-element group 946 branch  place  bypass 
    -- predecessors 945 
    -- successors 947 949 
    -- members (1) 
      -- 	branch_block_stmt_2042/R_orx_xcondx_xix_xi_3488_place
      -- 
    cp_elements(946) <= cp_elements(945);
    -- CP-element group 947 transition  bypass 
    -- predecessors 946 
    -- successors 948 
    -- members (1) 
      -- 	branch_block_stmt_2042/if_stmt_3487_if_link/$entry
      -- 
    cp_elements(947) <= cp_elements(946);
    -- CP-element group 948 transition  place  input  bypass 
    -- predecessors 947 
    -- successors 2172 
    -- members (3) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi_udiv32x_xexitx_xix_xi
      -- 	branch_block_stmt_2042/if_stmt_3487_if_link/$exit
      -- 	branch_block_stmt_2042/if_stmt_3487_if_link/if_choice_transition
      -- 
    if_choice_transition_14198_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_3487_branch_ack_1, ack => cp_elements(948)); -- 
    -- CP-element group 949 transition  bypass 
    -- predecessors 946 
    -- successors 950 
    -- members (1) 
      -- 	branch_block_stmt_2042/if_stmt_3487_else_link/$entry
      -- 
    cp_elements(949) <= cp_elements(946);
    -- CP-element group 950 transition  place  input  bypass 
    -- predecessors 949 
    -- successors 2215 
    -- members (3) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi_udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi
      -- 	branch_block_stmt_2042/if_stmt_3487_else_link/$exit
      -- 	branch_block_stmt_2042/if_stmt_3487_else_link/else_choice_transition
      -- 
    else_choice_transition_14202_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_3487_branch_ack_0, ack => cp_elements(950)); -- 
    -- CP-element group 951 fork  transition  bypass 
    -- predecessors 58 
    -- successors 952 953 957 958 962 963 
    -- members (1) 
      -- 	branch_block_stmt_2042/assign_stmt_3508_to_assign_stmt_3518/$entry
      -- 
    cp_elements(951) <= cp_elements(58);
    -- CP-element group 952 transition  output  bypass 
    -- predecessors 951 
    -- successors 955 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_3508_to_assign_stmt_3518/ADD_u32_u32_3507_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_3508_to_assign_stmt_3518/ADD_u32_u32_3507_Update/$entry
      -- 	branch_block_stmt_2042/assign_stmt_3508_to_assign_stmt_3518/ADD_u32_u32_3507_Update/cr
      -- 
    cp_elements(952) <= cp_elements(951);
    cr_14224_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(952), ack => ADD_u32_u32_3507_inst_req_1); -- 
    -- CP-element group 953 transition  output  bypass 
    -- predecessors 951 
    -- successors 954 
    -- members (7) 
      -- 	branch_block_stmt_2042/assign_stmt_3508_to_assign_stmt_3518/ADD_u32_u32_3507_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_3508_to_assign_stmt_3518/R_iNsTr_89_3504_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_3508_to_assign_stmt_3518/R_iNsTr_89_3504_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3508_to_assign_stmt_3518/R_iNsTr_89_3504_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_3508_to_assign_stmt_3518/R_iNsTr_89_3504_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3508_to_assign_stmt_3518/ADD_u32_u32_3507_Sample/$entry
      -- 	branch_block_stmt_2042/assign_stmt_3508_to_assign_stmt_3518/ADD_u32_u32_3507_Sample/rr
      -- 
    cp_elements(953) <= cp_elements(951);
    rr_14219_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(953), ack => ADD_u32_u32_3507_inst_req_0); -- 
    -- CP-element group 954 transition  input  bypass 
    -- predecessors 953 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_3508_to_assign_stmt_3518/ADD_u32_u32_3507_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3508_to_assign_stmt_3518/ADD_u32_u32_3507_Sample/$exit
      -- 	branch_block_stmt_2042/assign_stmt_3508_to_assign_stmt_3518/ADD_u32_u32_3507_Sample/ra
      -- 
    ra_14220_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u32_u32_3507_inst_ack_0, ack => cp_elements(954)); -- 
    -- CP-element group 955 transition  input  bypass 
    -- predecessors 952 
    -- successors 956 
    -- members (7) 
      -- 	branch_block_stmt_2042/assign_stmt_3508_to_assign_stmt_3518/ADD_u32_u32_3507_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3508_to_assign_stmt_3518/ADD_u32_u32_3507_Update/$exit
      -- 	branch_block_stmt_2042/assign_stmt_3508_to_assign_stmt_3518/ADD_u32_u32_3507_Update/ca
      -- 	branch_block_stmt_2042/assign_stmt_3508_to_assign_stmt_3518/R_tmp21x_xix_xi_3510_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_3508_to_assign_stmt_3518/R_tmp21x_xix_xi_3510_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3508_to_assign_stmt_3518/R_tmp21x_xix_xi_3510_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_3508_to_assign_stmt_3518/R_tmp21x_xix_xi_3510_update_completed_
      -- 
    ca_14225_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u32_u32_3507_inst_ack_1, ack => cp_elements(955)); -- 
    -- CP-element group 956 join  transition  output  bypass 
    -- predecessors 955 958 
    -- successors 959 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_3508_to_assign_stmt_3518/SUB_u32_u32_3512_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_3508_to_assign_stmt_3518/SUB_u32_u32_3512_Sample/$entry
      -- 	branch_block_stmt_2042/assign_stmt_3508_to_assign_stmt_3518/SUB_u32_u32_3512_Sample/rr
      -- 
    cp_element_group_956: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 20) := "cp_element_group_956"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(955) & cp_elements(958);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(956), clk => clk, reset => reset); --
    end block;
    rr_14241_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(956), ack => SUB_u32_u32_3512_inst_req_0); -- 
    -- CP-element group 957 transition  output  bypass 
    -- predecessors 951 
    -- successors 960 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_3508_to_assign_stmt_3518/SUB_u32_u32_3512_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_3508_to_assign_stmt_3518/SUB_u32_u32_3512_Update/$entry
      -- 	branch_block_stmt_2042/assign_stmt_3508_to_assign_stmt_3518/SUB_u32_u32_3512_Update/cr
      -- 
    cp_elements(957) <= cp_elements(951);
    cr_14246_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(957), ack => SUB_u32_u32_3512_inst_req_1); -- 
    -- CP-element group 958 transition  bypass 
    -- predecessors 951 
    -- successors 956 
    -- members (4) 
      -- 	branch_block_stmt_2042/assign_stmt_3508_to_assign_stmt_3518/R_iNsTr_91_3511_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_3508_to_assign_stmt_3518/R_iNsTr_91_3511_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3508_to_assign_stmt_3518/R_iNsTr_91_3511_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_3508_to_assign_stmt_3518/R_iNsTr_91_3511_update_completed_
      -- 
    cp_elements(958) <= cp_elements(951);
    -- CP-element group 959 transition  input  bypass 
    -- predecessors 956 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_3508_to_assign_stmt_3518/SUB_u32_u32_3512_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3508_to_assign_stmt_3518/SUB_u32_u32_3512_Sample/$exit
      -- 	branch_block_stmt_2042/assign_stmt_3508_to_assign_stmt_3518/SUB_u32_u32_3512_Sample/ra
      -- 
    ra_14242_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => SUB_u32_u32_3512_inst_ack_0, ack => cp_elements(959)); -- 
    -- CP-element group 960 transition  input  bypass 
    -- predecessors 957 
    -- successors 961 
    -- members (7) 
      -- 	branch_block_stmt_2042/assign_stmt_3508_to_assign_stmt_3518/SUB_u32_u32_3512_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3508_to_assign_stmt_3518/SUB_u32_u32_3512_Update/$exit
      -- 	branch_block_stmt_2042/assign_stmt_3508_to_assign_stmt_3518/SUB_u32_u32_3512_Update/ca
      -- 	branch_block_stmt_2042/assign_stmt_3508_to_assign_stmt_3518/R_tmp25x_xix_xi_3515_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_3508_to_assign_stmt_3518/R_tmp25x_xix_xi_3515_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3508_to_assign_stmt_3518/R_tmp25x_xix_xi_3515_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_3508_to_assign_stmt_3518/R_tmp25x_xix_xi_3515_update_completed_
      -- 
    ca_14247_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => SUB_u32_u32_3512_inst_ack_1, ack => cp_elements(960)); -- 
    -- CP-element group 961 join  transition  output  bypass 
    -- predecessors 960 963 
    -- successors 964 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_3508_to_assign_stmt_3518/SUB_u32_u32_3517_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_3508_to_assign_stmt_3518/SUB_u32_u32_3517_Sample/$entry
      -- 	branch_block_stmt_2042/assign_stmt_3508_to_assign_stmt_3518/SUB_u32_u32_3517_Sample/rr
      -- 
    cp_element_group_961: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 20) := "cp_element_group_961"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(960) & cp_elements(963);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(961), clk => clk, reset => reset); --
    end block;
    rr_14263_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(961), ack => SUB_u32_u32_3517_inst_req_0); -- 
    -- CP-element group 962 transition  output  bypass 
    -- predecessors 951 
    -- successors 965 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_3508_to_assign_stmt_3518/SUB_u32_u32_3517_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_3508_to_assign_stmt_3518/SUB_u32_u32_3517_Update/$entry
      -- 	branch_block_stmt_2042/assign_stmt_3508_to_assign_stmt_3518/SUB_u32_u32_3517_Update/cr
      -- 
    cp_elements(962) <= cp_elements(951);
    cr_14268_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(962), ack => SUB_u32_u32_3517_inst_req_1); -- 
    -- CP-element group 963 transition  bypass 
    -- predecessors 951 
    -- successors 961 
    -- members (4) 
      -- 	branch_block_stmt_2042/assign_stmt_3508_to_assign_stmt_3518/R_xx_xlcssa5_3516_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_3508_to_assign_stmt_3518/R_xx_xlcssa5_3516_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3508_to_assign_stmt_3518/R_xx_xlcssa5_3516_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_3508_to_assign_stmt_3518/R_xx_xlcssa5_3516_update_completed_
      -- 
    cp_elements(963) <= cp_elements(951);
    -- CP-element group 964 transition  input  bypass 
    -- predecessors 961 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_3508_to_assign_stmt_3518/SUB_u32_u32_3517_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3508_to_assign_stmt_3518/SUB_u32_u32_3517_Sample/$exit
      -- 	branch_block_stmt_2042/assign_stmt_3508_to_assign_stmt_3518/SUB_u32_u32_3517_Sample/ra
      -- 
    ra_14264_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => SUB_u32_u32_3517_inst_ack_0, ack => cp_elements(964)); -- 
    -- CP-element group 965 transition  place  input  bypass 
    -- predecessors 962 
    -- successors 2260 
    -- members (6) 
      -- 	branch_block_stmt_2042/assign_stmt_3508_to_assign_stmt_3518__exit__
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi_xx_xcritedgex_xix_xi
      -- 	branch_block_stmt_2042/assign_stmt_3508_to_assign_stmt_3518/$exit
      -- 	branch_block_stmt_2042/assign_stmt_3508_to_assign_stmt_3518/SUB_u32_u32_3517_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3508_to_assign_stmt_3518/SUB_u32_u32_3517_Update/$exit
      -- 	branch_block_stmt_2042/assign_stmt_3508_to_assign_stmt_3518/SUB_u32_u32_3517_Update/ca
      -- 
    ca_14269_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => SUB_u32_u32_3517_inst_ack_1, ack => cp_elements(965)); -- 
    -- CP-element group 966 fork  transition  bypass 
    -- predecessors 59 
    -- successors 967 968 971 972 975 979 980 984 987 
    -- members (1) 
      -- 	branch_block_stmt_2042/assign_stmt_3539_to_assign_stmt_3565/$entry
      -- 
    cp_elements(966) <= cp_elements(59);
    -- CP-element group 967 transition  output  bypass 
    -- predecessors 966 
    -- successors 970 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_3539_to_assign_stmt_3565/AND_u32_u32_3538_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_3539_to_assign_stmt_3565/AND_u32_u32_3538_Update/$entry
      -- 	branch_block_stmt_2042/assign_stmt_3539_to_assign_stmt_3565/AND_u32_u32_3538_Update/cr
      -- 
    cp_elements(967) <= cp_elements(966);
    cr_14289_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(967), ack => AND_u32_u32_3538_inst_req_1); -- 
    -- CP-element group 968 transition  output  bypass 
    -- predecessors 966 
    -- successors 969 
    -- members (7) 
      -- 	branch_block_stmt_2042/assign_stmt_3539_to_assign_stmt_3565/AND_u32_u32_3538_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_3539_to_assign_stmt_3565/R_tempx_x0x_xlcssax_xix_xi_3535_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_3539_to_assign_stmt_3565/R_tempx_x0x_xlcssax_xix_xi_3535_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3539_to_assign_stmt_3565/R_tempx_x0x_xlcssax_xix_xi_3535_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_3539_to_assign_stmt_3565/R_tempx_x0x_xlcssax_xix_xi_3535_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3539_to_assign_stmt_3565/AND_u32_u32_3538_Sample/$entry
      -- 	branch_block_stmt_2042/assign_stmt_3539_to_assign_stmt_3565/AND_u32_u32_3538_Sample/rr
      -- 
    cp_elements(968) <= cp_elements(966);
    rr_14284_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(968), ack => AND_u32_u32_3538_inst_req_0); -- 
    -- CP-element group 969 transition  input  bypass 
    -- predecessors 968 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_3539_to_assign_stmt_3565/AND_u32_u32_3538_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3539_to_assign_stmt_3565/AND_u32_u32_3538_Sample/$exit
      -- 	branch_block_stmt_2042/assign_stmt_3539_to_assign_stmt_3565/AND_u32_u32_3538_Sample/ra
      -- 
    ra_14285_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => AND_u32_u32_3538_inst_ack_0, ack => cp_elements(969)); -- 
    -- CP-element group 970 transition  input  bypass 
    -- predecessors 967 
    -- successors 978 
    -- members (7) 
      -- 	branch_block_stmt_2042/assign_stmt_3539_to_assign_stmt_3565/AND_u32_u32_3538_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3539_to_assign_stmt_3565/AND_u32_u32_3538_Update/$exit
      -- 	branch_block_stmt_2042/assign_stmt_3539_to_assign_stmt_3565/AND_u32_u32_3538_Update/ca
      -- 	branch_block_stmt_2042/assign_stmt_3539_to_assign_stmt_3565/R_iNsTr_158_3553_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_3539_to_assign_stmt_3565/R_iNsTr_158_3553_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3539_to_assign_stmt_3565/R_iNsTr_158_3553_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_3539_to_assign_stmt_3565/R_iNsTr_158_3553_update_completed_
      -- 
    ca_14290_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => AND_u32_u32_3538_inst_ack_1, ack => cp_elements(970)); -- 
    -- CP-element group 971 transition  output  bypass 
    -- predecessors 966 
    -- successors 974 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_3539_to_assign_stmt_3565/SHL_u32_u32_3544_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_3539_to_assign_stmt_3565/SHL_u32_u32_3544_Update/$entry
      -- 	branch_block_stmt_2042/assign_stmt_3539_to_assign_stmt_3565/SHL_u32_u32_3544_Update/cr
      -- 
    cp_elements(971) <= cp_elements(966);
    cr_14307_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(971), ack => SHL_u32_u32_3544_inst_req_1); -- 
    -- CP-element group 972 transition  output  bypass 
    -- predecessors 966 
    -- successors 973 
    -- members (7) 
      -- 	branch_block_stmt_2042/assign_stmt_3539_to_assign_stmt_3565/SHL_u32_u32_3544_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_3539_to_assign_stmt_3565/R_expx_x0x_xlcssax_xix_xi_3541_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_3539_to_assign_stmt_3565/R_expx_x0x_xlcssax_xix_xi_3541_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3539_to_assign_stmt_3565/R_expx_x0x_xlcssax_xix_xi_3541_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_3539_to_assign_stmt_3565/R_expx_x0x_xlcssax_xix_xi_3541_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3539_to_assign_stmt_3565/SHL_u32_u32_3544_Sample/$entry
      -- 	branch_block_stmt_2042/assign_stmt_3539_to_assign_stmt_3565/SHL_u32_u32_3544_Sample/rr
      -- 
    cp_elements(972) <= cp_elements(966);
    rr_14302_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(972), ack => SHL_u32_u32_3544_inst_req_0); -- 
    -- CP-element group 973 transition  input  bypass 
    -- predecessors 972 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_3539_to_assign_stmt_3565/SHL_u32_u32_3544_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3539_to_assign_stmt_3565/SHL_u32_u32_3544_Sample/$exit
      -- 	branch_block_stmt_2042/assign_stmt_3539_to_assign_stmt_3565/SHL_u32_u32_3544_Sample/ra
      -- 
    ra_14303_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => SHL_u32_u32_3544_inst_ack_0, ack => cp_elements(973)); -- 
    -- CP-element group 974 transition  input  output  bypass 
    -- predecessors 971 
    -- successors 976 
    -- members (10) 
      -- 	branch_block_stmt_2042/assign_stmt_3539_to_assign_stmt_3565/SHL_u32_u32_3544_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3539_to_assign_stmt_3565/SHL_u32_u32_3544_Update/$exit
      -- 	branch_block_stmt_2042/assign_stmt_3539_to_assign_stmt_3565/SHL_u32_u32_3544_Update/ca
      -- 	branch_block_stmt_2042/assign_stmt_3539_to_assign_stmt_3565/ADD_u32_u32_3550_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_3539_to_assign_stmt_3565/R_iNsTr_159_3547_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_3539_to_assign_stmt_3565/R_iNsTr_159_3547_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3539_to_assign_stmt_3565/R_iNsTr_159_3547_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_3539_to_assign_stmt_3565/R_iNsTr_159_3547_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3539_to_assign_stmt_3565/ADD_u32_u32_3550_Sample/$entry
      -- 	branch_block_stmt_2042/assign_stmt_3539_to_assign_stmt_3565/ADD_u32_u32_3550_Sample/rr
      -- 
    ca_14308_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => SHL_u32_u32_3544_inst_ack_1, ack => cp_elements(974)); -- 
    rr_14320_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(974), ack => ADD_u32_u32_3550_inst_req_0); -- 
    -- CP-element group 975 transition  output  bypass 
    -- predecessors 966 
    -- successors 977 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_3539_to_assign_stmt_3565/ADD_u32_u32_3550_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_3539_to_assign_stmt_3565/ADD_u32_u32_3550_Update/$entry
      -- 	branch_block_stmt_2042/assign_stmt_3539_to_assign_stmt_3565/ADD_u32_u32_3550_Update/cr
      -- 
    cp_elements(975) <= cp_elements(966);
    cr_14325_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(975), ack => ADD_u32_u32_3550_inst_req_1); -- 
    -- CP-element group 976 transition  input  bypass 
    -- predecessors 974 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_3539_to_assign_stmt_3565/ADD_u32_u32_3550_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3539_to_assign_stmt_3565/ADD_u32_u32_3550_Sample/$exit
      -- 	branch_block_stmt_2042/assign_stmt_3539_to_assign_stmt_3565/ADD_u32_u32_3550_Sample/ra
      -- 
    ra_14321_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u32_u32_3550_inst_ack_0, ack => cp_elements(976)); -- 
    -- CP-element group 977 transition  input  bypass 
    -- predecessors 975 
    -- successors 983 
    -- members (7) 
      -- 	branch_block_stmt_2042/assign_stmt_3539_to_assign_stmt_3565/ADD_u32_u32_3550_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3539_to_assign_stmt_3565/ADD_u32_u32_3550_Update/$exit
      -- 	branch_block_stmt_2042/assign_stmt_3539_to_assign_stmt_3565/ADD_u32_u32_3550_Update/ca
      -- 	branch_block_stmt_2042/assign_stmt_3539_to_assign_stmt_3565/R_iNsTr_160_3559_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_3539_to_assign_stmt_3565/R_iNsTr_160_3559_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3539_to_assign_stmt_3565/R_iNsTr_160_3559_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_3539_to_assign_stmt_3565/R_iNsTr_160_3559_update_completed_
      -- 
    ca_14326_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u32_u32_3550_inst_ack_1, ack => cp_elements(977)); -- 
    -- CP-element group 978 join  transition  output  bypass 
    -- predecessors 970 980 
    -- successors 981 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_3539_to_assign_stmt_3565/OR_u32_u32_3555_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_3539_to_assign_stmt_3565/OR_u32_u32_3555_Sample/$entry
      -- 	branch_block_stmt_2042/assign_stmt_3539_to_assign_stmt_3565/OR_u32_u32_3555_Sample/rr
      -- 
    cp_element_group_978: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 20) := "cp_element_group_978"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(970) & cp_elements(980);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(978), clk => clk, reset => reset); --
    end block;
    rr_14342_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(978), ack => OR_u32_u32_3555_inst_req_0); -- 
    -- CP-element group 979 transition  output  bypass 
    -- predecessors 966 
    -- successors 982 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_3539_to_assign_stmt_3565/OR_u32_u32_3555_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_3539_to_assign_stmt_3565/OR_u32_u32_3555_Update/$entry
      -- 	branch_block_stmt_2042/assign_stmt_3539_to_assign_stmt_3565/OR_u32_u32_3555_Update/cr
      -- 
    cp_elements(979) <= cp_elements(966);
    cr_14347_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(979), ack => OR_u32_u32_3555_inst_req_1); -- 
    -- CP-element group 980 transition  bypass 
    -- predecessors 966 
    -- successors 978 
    -- members (4) 
      -- 	branch_block_stmt_2042/assign_stmt_3539_to_assign_stmt_3565/R_iNsTr_99_3554_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_3539_to_assign_stmt_3565/R_iNsTr_99_3554_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3539_to_assign_stmt_3565/R_iNsTr_99_3554_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_3539_to_assign_stmt_3565/R_iNsTr_99_3554_update_completed_
      -- 
    cp_elements(980) <= cp_elements(966);
    -- CP-element group 981 transition  input  bypass 
    -- predecessors 978 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_3539_to_assign_stmt_3565/OR_u32_u32_3555_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3539_to_assign_stmt_3565/OR_u32_u32_3555_Sample/$exit
      -- 	branch_block_stmt_2042/assign_stmt_3539_to_assign_stmt_3565/OR_u32_u32_3555_Sample/ra
      -- 
    ra_14343_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => OR_u32_u32_3555_inst_ack_0, ack => cp_elements(981)); -- 
    -- CP-element group 982 transition  input  bypass 
    -- predecessors 979 
    -- successors 983 
    -- members (7) 
      -- 	branch_block_stmt_2042/assign_stmt_3539_to_assign_stmt_3565/OR_u32_u32_3555_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3539_to_assign_stmt_3565/OR_u32_u32_3555_Update/$exit
      -- 	branch_block_stmt_2042/assign_stmt_3539_to_assign_stmt_3565/OR_u32_u32_3555_Update/ca
      -- 	branch_block_stmt_2042/assign_stmt_3539_to_assign_stmt_3565/R_iNsTr_161_3558_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_3539_to_assign_stmt_3565/R_iNsTr_161_3558_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3539_to_assign_stmt_3565/R_iNsTr_161_3558_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_3539_to_assign_stmt_3565/R_iNsTr_161_3558_update_completed_
      -- 
    ca_14348_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => OR_u32_u32_3555_inst_ack_1, ack => cp_elements(982)); -- 
    -- CP-element group 983 join  transition  output  bypass 
    -- predecessors 977 982 
    -- successors 985 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_3539_to_assign_stmt_3565/OR_u32_u32_3560_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_3539_to_assign_stmt_3565/OR_u32_u32_3560_Sample/$entry
      -- 	branch_block_stmt_2042/assign_stmt_3539_to_assign_stmt_3565/OR_u32_u32_3560_Sample/rr
      -- 
    cp_element_group_983: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 20) := "cp_element_group_983"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(977) & cp_elements(982);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(983), clk => clk, reset => reset); --
    end block;
    rr_14364_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(983), ack => OR_u32_u32_3560_inst_req_0); -- 
    -- CP-element group 984 transition  output  bypass 
    -- predecessors 966 
    -- successors 986 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_3539_to_assign_stmt_3565/OR_u32_u32_3560_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_3539_to_assign_stmt_3565/OR_u32_u32_3560_Update/$entry
      -- 	branch_block_stmt_2042/assign_stmt_3539_to_assign_stmt_3565/OR_u32_u32_3560_Update/cr
      -- 
    cp_elements(984) <= cp_elements(966);
    cr_14369_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(984), ack => OR_u32_u32_3560_inst_req_1); -- 
    -- CP-element group 985 transition  input  bypass 
    -- predecessors 983 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_3539_to_assign_stmt_3565/OR_u32_u32_3560_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3539_to_assign_stmt_3565/OR_u32_u32_3560_Sample/$exit
      -- 	branch_block_stmt_2042/assign_stmt_3539_to_assign_stmt_3565/OR_u32_u32_3560_Sample/ra
      -- 
    ra_14365_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => OR_u32_u32_3560_inst_ack_0, ack => cp_elements(985)); -- 
    -- CP-element group 986 transition  input  output  bypass 
    -- predecessors 984 
    -- successors 988 
    -- members (10) 
      -- 	branch_block_stmt_2042/assign_stmt_3539_to_assign_stmt_3565/R_iNsTr_162_3563_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3539_to_assign_stmt_3565/OR_u32_u32_3560_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3539_to_assign_stmt_3565/OR_u32_u32_3560_Update/$exit
      -- 	branch_block_stmt_2042/assign_stmt_3539_to_assign_stmt_3565/OR_u32_u32_3560_Update/ca
      -- 	branch_block_stmt_2042/assign_stmt_3539_to_assign_stmt_3565/type_cast_3564_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_3539_to_assign_stmt_3565/R_iNsTr_162_3563_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_3539_to_assign_stmt_3565/R_iNsTr_162_3563_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3539_to_assign_stmt_3565/R_iNsTr_162_3563_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_3539_to_assign_stmt_3565/type_cast_3564_Sample/$entry
      -- 	branch_block_stmt_2042/assign_stmt_3539_to_assign_stmt_3565/type_cast_3564_Sample/rr
      -- 
    ca_14370_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => OR_u32_u32_3560_inst_ack_1, ack => cp_elements(986)); -- 
    rr_14382_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(986), ack => type_cast_3564_inst_req_0); -- 
    -- CP-element group 987 transition  output  bypass 
    -- predecessors 966 
    -- successors 989 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_3539_to_assign_stmt_3565/type_cast_3564_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_3539_to_assign_stmt_3565/type_cast_3564_Update/$entry
      -- 	branch_block_stmt_2042/assign_stmt_3539_to_assign_stmt_3565/type_cast_3564_Update/cr
      -- 
    cp_elements(987) <= cp_elements(966);
    cr_14387_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(987), ack => type_cast_3564_inst_req_1); -- 
    -- CP-element group 988 transition  input  bypass 
    -- predecessors 986 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_3539_to_assign_stmt_3565/type_cast_3564_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3539_to_assign_stmt_3565/type_cast_3564_Sample/$exit
      -- 	branch_block_stmt_2042/assign_stmt_3539_to_assign_stmt_3565/type_cast_3564_Sample/ra
      -- 
    ra_14383_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3564_inst_ack_0, ack => cp_elements(988)); -- 
    -- CP-element group 989 fork  transition  place  input  bypass 
    -- predecessors 987 
    -- successors 2294 2296 
    -- members (11) 
      -- 	branch_block_stmt_2042/assign_stmt_3539_to_assign_stmt_3565__exit__
      -- 	branch_block_stmt_2042/xx_xcritedgex_xix_xi_iq_err_calcx_xexit
      -- 	branch_block_stmt_2042/assign_stmt_3539_to_assign_stmt_3565/$exit
      -- 	branch_block_stmt_2042/assign_stmt_3539_to_assign_stmt_3565/type_cast_3564_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3539_to_assign_stmt_3565/type_cast_3564_Update/$exit
      -- 	branch_block_stmt_2042/assign_stmt_3539_to_assign_stmt_3565/type_cast_3564_Update/ca
      -- 	branch_block_stmt_2042/xx_xcritedgex_xix_xi_iq_err_calcx_xexit_PhiReq/$entry
      -- 	branch_block_stmt_2042/xx_xcritedgex_xix_xi_iq_err_calcx_xexit_PhiReq/phi_stmt_3568/$entry
      -- 	branch_block_stmt_2042/xx_xcritedgex_xix_xi_iq_err_calcx_xexit_PhiReq/phi_stmt_3568/phi_stmt_3568_sources/$entry
      -- 	branch_block_stmt_2042/xx_xcritedgex_xix_xi_iq_err_calcx_xexit_PhiReq/phi_stmt_3568/phi_stmt_3568_sources/type_cast_3571/$entry
      -- 	branch_block_stmt_2042/xx_xcritedgex_xix_xi_iq_err_calcx_xexit_PhiReq/phi_stmt_3568/phi_stmt_3568_sources/type_cast_3571/SplitProtocol/$entry
      -- 
    ca_14388_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3564_inst_ack_1, ack => cp_elements(989)); -- 
    -- CP-element group 990 fork  transition  bypass 
    -- predecessors 2301 
    -- successors 992 993 994 997 1001 1002 1005 1008 
    -- members (1) 
      -- 	branch_block_stmt_2042/assign_stmt_3580_to_assign_stmt_3603/$entry
      -- 
    cp_elements(990) <= cp_elements(2301);
    -- CP-element group 991 join  transition  output  bypass 
    -- predecessors 993 994 
    -- successors 995 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_3580_to_assign_stmt_3603/SUB_f32_f32_3579_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_3580_to_assign_stmt_3603/SUB_f32_f32_3579_Sample/$entry
      -- 	branch_block_stmt_2042/assign_stmt_3580_to_assign_stmt_3603/SUB_f32_f32_3579_Sample/rr
      -- 
    cp_element_group_991: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 20) := "cp_element_group_991"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(993) & cp_elements(994);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(991), clk => clk, reset => reset); --
    end block;
    rr_14407_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(991), ack => SUB_f32_f32_3579_inst_req_0); -- 
    -- CP-element group 992 transition  output  bypass 
    -- predecessors 990 
    -- successors 996 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_3580_to_assign_stmt_3603/SUB_f32_f32_3579_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_3580_to_assign_stmt_3603/SUB_f32_f32_3579_Update/$entry
      -- 	branch_block_stmt_2042/assign_stmt_3580_to_assign_stmt_3603/SUB_f32_f32_3579_Update/cr
      -- 
    cp_elements(992) <= cp_elements(990);
    cr_14412_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(992), ack => SUB_f32_f32_3579_inst_req_1); -- 
    -- CP-element group 993 transition  bypass 
    -- predecessors 990 
    -- successors 991 
    -- members (4) 
      -- 	branch_block_stmt_2042/assign_stmt_3580_to_assign_stmt_3603/R_flux_refx_x0_3577_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_3580_to_assign_stmt_3603/R_flux_refx_x0_3577_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3580_to_assign_stmt_3603/R_flux_refx_x0_3577_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_3580_to_assign_stmt_3603/R_flux_refx_x0_3577_update_completed_
      -- 
    cp_elements(993) <= cp_elements(990);
    -- CP-element group 994 transition  bypass 
    -- predecessors 990 
    -- successors 991 
    -- members (4) 
      -- 	branch_block_stmt_2042/assign_stmt_3580_to_assign_stmt_3603/R_iNsTr_42_3578_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_3580_to_assign_stmt_3603/R_iNsTr_42_3578_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3580_to_assign_stmt_3603/R_iNsTr_42_3578_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_3580_to_assign_stmt_3603/R_iNsTr_42_3578_update_completed_
      -- 
    cp_elements(994) <= cp_elements(990);
    -- CP-element group 995 transition  input  bypass 
    -- predecessors 991 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_3580_to_assign_stmt_3603/SUB_f32_f32_3579_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3580_to_assign_stmt_3603/SUB_f32_f32_3579_Sample/$exit
      -- 	branch_block_stmt_2042/assign_stmt_3580_to_assign_stmt_3603/SUB_f32_f32_3579_Sample/ra
      -- 
    ra_14408_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => SUB_f32_f32_3579_inst_ack_0, ack => cp_elements(995)); -- 
    -- CP-element group 996 transition  input  output  bypass 
    -- predecessors 992 
    -- successors 998 
    -- members (10) 
      -- 	branch_block_stmt_2042/assign_stmt_3580_to_assign_stmt_3603/SUB_f32_f32_3579_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3580_to_assign_stmt_3603/SUB_f32_f32_3579_Update/$exit
      -- 	branch_block_stmt_2042/assign_stmt_3580_to_assign_stmt_3603/SUB_f32_f32_3579_Update/ca
      -- 	branch_block_stmt_2042/assign_stmt_3580_to_assign_stmt_3603/MUL_f32_f32_3585_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_3580_to_assign_stmt_3603/R_iNsTr_82_3582_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_3580_to_assign_stmt_3603/R_iNsTr_82_3582_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3580_to_assign_stmt_3603/R_iNsTr_82_3582_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_3580_to_assign_stmt_3603/R_iNsTr_82_3582_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3580_to_assign_stmt_3603/MUL_f32_f32_3585_Sample/$entry
      -- 	branch_block_stmt_2042/assign_stmt_3580_to_assign_stmt_3603/MUL_f32_f32_3585_Sample/rr
      -- 
    ca_14413_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => SUB_f32_f32_3579_inst_ack_1, ack => cp_elements(996)); -- 
    rr_14425_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(996), ack => MUL_f32_f32_3585_inst_req_0); -- 
    -- CP-element group 997 transition  output  bypass 
    -- predecessors 990 
    -- successors 999 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_3580_to_assign_stmt_3603/MUL_f32_f32_3585_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_3580_to_assign_stmt_3603/MUL_f32_f32_3585_Update/$entry
      -- 	branch_block_stmt_2042/assign_stmt_3580_to_assign_stmt_3603/MUL_f32_f32_3585_Update/cr
      -- 
    cp_elements(997) <= cp_elements(990);
    cr_14430_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(997), ack => MUL_f32_f32_3585_inst_req_1); -- 
    -- CP-element group 998 transition  input  bypass 
    -- predecessors 996 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_3580_to_assign_stmt_3603/MUL_f32_f32_3585_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3580_to_assign_stmt_3603/MUL_f32_f32_3585_Sample/$exit
      -- 	branch_block_stmt_2042/assign_stmt_3580_to_assign_stmt_3603/MUL_f32_f32_3585_Sample/ra
      -- 
    ra_14426_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => MUL_f32_f32_3585_inst_ack_0, ack => cp_elements(998)); -- 
    -- CP-element group 999 transition  input  bypass 
    -- predecessors 997 
    -- successors 1000 
    -- members (7) 
      -- 	branch_block_stmt_2042/assign_stmt_3580_to_assign_stmt_3603/MUL_f32_f32_3585_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3580_to_assign_stmt_3603/MUL_f32_f32_3585_Update/$exit
      -- 	branch_block_stmt_2042/assign_stmt_3580_to_assign_stmt_3603/MUL_f32_f32_3585_Update/ca
      -- 	branch_block_stmt_2042/assign_stmt_3580_to_assign_stmt_3603/R_iNsTr_83_3588_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_3580_to_assign_stmt_3603/R_iNsTr_83_3588_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3580_to_assign_stmt_3603/R_iNsTr_83_3588_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_3580_to_assign_stmt_3603/R_iNsTr_83_3588_update_completed_
      -- 
    ca_14431_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => MUL_f32_f32_3585_inst_ack_1, ack => cp_elements(999)); -- 
    -- CP-element group 1000 join  transition  output  bypass 
    -- predecessors 999 1002 
    -- successors 1003 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_3580_to_assign_stmt_3603/ADD_f32_f32_3590_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_3580_to_assign_stmt_3603/ADD_f32_f32_3590_Sample/$entry
      -- 	branch_block_stmt_2042/assign_stmt_3580_to_assign_stmt_3603/ADD_f32_f32_3590_Sample/rr
      -- 
    cp_element_group_1000: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1000"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(999) & cp_elements(1002);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1000), clk => clk, reset => reset); --
    end block;
    rr_14447_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1000), ack => ADD_f32_f32_3590_inst_req_0); -- 
    -- CP-element group 1001 transition  output  bypass 
    -- predecessors 990 
    -- successors 1004 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_3580_to_assign_stmt_3603/ADD_f32_f32_3590_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_3580_to_assign_stmt_3603/ADD_f32_f32_3590_Update/$entry
      -- 	branch_block_stmt_2042/assign_stmt_3580_to_assign_stmt_3603/ADD_f32_f32_3590_Update/cr
      -- 
    cp_elements(1001) <= cp_elements(990);
    cr_14452_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1001), ack => ADD_f32_f32_3590_inst_req_1); -- 
    -- CP-element group 1002 transition  bypass 
    -- predecessors 990 
    -- successors 1000 
    -- members (4) 
      -- 	branch_block_stmt_2042/assign_stmt_3580_to_assign_stmt_3603/R_int_flux_errx_x0_3589_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_3580_to_assign_stmt_3603/R_int_flux_errx_x0_3589_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3580_to_assign_stmt_3603/R_int_flux_errx_x0_3589_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_3580_to_assign_stmt_3603/R_int_flux_errx_x0_3589_update_completed_
      -- 
    cp_elements(1002) <= cp_elements(990);
    -- CP-element group 1003 transition  input  bypass 
    -- predecessors 1000 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_3580_to_assign_stmt_3603/ADD_f32_f32_3590_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3580_to_assign_stmt_3603/ADD_f32_f32_3590_Sample/$exit
      -- 	branch_block_stmt_2042/assign_stmt_3580_to_assign_stmt_3603/ADD_f32_f32_3590_Sample/ra
      -- 
    ra_14448_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_f32_f32_3590_inst_ack_0, ack => cp_elements(1003)); -- 
    -- CP-element group 1004 transition  input  output  bypass 
    -- predecessors 1001 
    -- successors 1006 
    -- members (10) 
      -- 	branch_block_stmt_2042/assign_stmt_3580_to_assign_stmt_3603/ADD_f32_f32_3590_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3580_to_assign_stmt_3603/ADD_f32_f32_3590_Update/$exit
      -- 	branch_block_stmt_2042/assign_stmt_3580_to_assign_stmt_3603/ADD_f32_f32_3590_Update/ca
      -- 	branch_block_stmt_2042/assign_stmt_3580_to_assign_stmt_3603/MUL_f32_f32_3596_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_3580_to_assign_stmt_3603/R_iNsTr_84_3593_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_3580_to_assign_stmt_3603/R_iNsTr_84_3593_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3580_to_assign_stmt_3603/R_iNsTr_84_3593_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_3580_to_assign_stmt_3603/R_iNsTr_84_3593_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3580_to_assign_stmt_3603/MUL_f32_f32_3596_Sample/$entry
      -- 	branch_block_stmt_2042/assign_stmt_3580_to_assign_stmt_3603/MUL_f32_f32_3596_Sample/rr
      -- 
    ca_14453_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_f32_f32_3590_inst_ack_1, ack => cp_elements(1004)); -- 
    rr_14465_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1004), ack => MUL_f32_f32_3596_inst_req_0); -- 
    -- CP-element group 1005 transition  output  bypass 
    -- predecessors 990 
    -- successors 1007 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_3580_to_assign_stmt_3603/MUL_f32_f32_3596_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_3580_to_assign_stmt_3603/MUL_f32_f32_3596_Update/$entry
      -- 	branch_block_stmt_2042/assign_stmt_3580_to_assign_stmt_3603/MUL_f32_f32_3596_Update/cr
      -- 
    cp_elements(1005) <= cp_elements(990);
    cr_14470_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1005), ack => MUL_f32_f32_3596_inst_req_1); -- 
    -- CP-element group 1006 transition  input  bypass 
    -- predecessors 1004 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_3580_to_assign_stmt_3603/MUL_f32_f32_3596_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3580_to_assign_stmt_3603/MUL_f32_f32_3596_Sample/$exit
      -- 	branch_block_stmt_2042/assign_stmt_3580_to_assign_stmt_3603/MUL_f32_f32_3596_Sample/ra
      -- 
    ra_14466_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => MUL_f32_f32_3596_inst_ack_0, ack => cp_elements(1006)); -- 
    -- CP-element group 1007 transition  input  output  bypass 
    -- predecessors 1005 
    -- successors 1009 
    -- members (10) 
      -- 	branch_block_stmt_2042/assign_stmt_3580_to_assign_stmt_3603/MUL_f32_f32_3596_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3580_to_assign_stmt_3603/MUL_f32_f32_3596_Update/$exit
      -- 	branch_block_stmt_2042/assign_stmt_3580_to_assign_stmt_3603/MUL_f32_f32_3596_Update/ca
      -- 	branch_block_stmt_2042/assign_stmt_3580_to_assign_stmt_3603/SLT_f32_u1_3602_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_3580_to_assign_stmt_3603/R_iNsTr_85_3599_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_3580_to_assign_stmt_3603/R_iNsTr_85_3599_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3580_to_assign_stmt_3603/R_iNsTr_85_3599_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_3580_to_assign_stmt_3603/R_iNsTr_85_3599_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3580_to_assign_stmt_3603/SLT_f32_u1_3602_Sample/$entry
      -- 	branch_block_stmt_2042/assign_stmt_3580_to_assign_stmt_3603/SLT_f32_u1_3602_Sample/rr
      -- 
    ca_14471_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => MUL_f32_f32_3596_inst_ack_1, ack => cp_elements(1007)); -- 
    rr_14483_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1007), ack => SLT_f32_u1_3602_inst_req_0); -- 
    -- CP-element group 1008 transition  output  bypass 
    -- predecessors 990 
    -- successors 1010 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_3580_to_assign_stmt_3603/SLT_f32_u1_3602_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_3580_to_assign_stmt_3603/SLT_f32_u1_3602_Update/$entry
      -- 	branch_block_stmt_2042/assign_stmt_3580_to_assign_stmt_3603/SLT_f32_u1_3602_Update/cr
      -- 
    cp_elements(1008) <= cp_elements(990);
    cr_14488_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1008), ack => SLT_f32_u1_3602_inst_req_1); -- 
    -- CP-element group 1009 transition  input  bypass 
    -- predecessors 1007 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_3580_to_assign_stmt_3603/SLT_f32_u1_3602_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3580_to_assign_stmt_3603/SLT_f32_u1_3602_Sample/$exit
      -- 	branch_block_stmt_2042/assign_stmt_3580_to_assign_stmt_3603/SLT_f32_u1_3602_Sample/ra
      -- 
    ra_14484_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => SLT_f32_u1_3602_inst_ack_0, ack => cp_elements(1009)); -- 
    -- CP-element group 1010 branch  transition  place  input  bypass 
    -- predecessors 1008 
    -- successors 1011 1012 
    -- members (6) 
      -- 	branch_block_stmt_2042/if_stmt_3604__entry__
      -- 	branch_block_stmt_2042/assign_stmt_3580_to_assign_stmt_3603__exit__
      -- 	branch_block_stmt_2042/assign_stmt_3580_to_assign_stmt_3603/$exit
      -- 	branch_block_stmt_2042/assign_stmt_3580_to_assign_stmt_3603/SLT_f32_u1_3602_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3580_to_assign_stmt_3603/SLT_f32_u1_3602_Update/$exit
      -- 	branch_block_stmt_2042/assign_stmt_3580_to_assign_stmt_3603/SLT_f32_u1_3602_Update/ca
      -- 
    ca_14489_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => SLT_f32_u1_3602_inst_ack_1, ack => cp_elements(1010)); -- 
    -- CP-element group 1011 transition  place  dead  bypass 
    -- predecessors 1010 
    -- successors 60 
    -- members (8) 
      -- 	branch_block_stmt_2042/merge_stmt_3610__entry__
      -- 	branch_block_stmt_2042/if_stmt_3604__exit__
      -- 	branch_block_stmt_2042/if_stmt_3604_dead_link/$entry
      -- 	branch_block_stmt_2042/if_stmt_3604_dead_link/$exit
      -- 	branch_block_stmt_2042/if_stmt_3604_dead_link/dead_transition
      -- 	branch_block_stmt_2042/merge_stmt_3610_dead_link/$entry
      -- 	branch_block_stmt_2042/merge_stmt_3610_dead_link/$exit
      -- 	branch_block_stmt_2042/merge_stmt_3610_dead_link/dead_transition
      -- 
    cp_elements(1011) <= false;
    -- CP-element group 1012 transition  output  bypass 
    -- predecessors 1010 
    -- successors 1013 
    -- members (3) 
      -- 	branch_block_stmt_2042/if_stmt_3604_eval_test/$entry
      -- 	branch_block_stmt_2042/if_stmt_3604_eval_test/$exit
      -- 	branch_block_stmt_2042/if_stmt_3604_eval_test/branch_req
      -- 
    cp_elements(1012) <= cp_elements(1010);
    branch_req_14497_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1012), ack => if_stmt_3604_branch_req_0); -- 
    -- CP-element group 1013 branch  place  bypass 
    -- predecessors 1012 
    -- successors 1014 1016 
    -- members (1) 
      -- 	branch_block_stmt_2042/R_iNsTr_86_3605_place
      -- 
    cp_elements(1013) <= cp_elements(1012);
    -- CP-element group 1014 transition  bypass 
    -- predecessors 1013 
    -- successors 1015 
    -- members (1) 
      -- 	branch_block_stmt_2042/if_stmt_3604_if_link/$entry
      -- 
    cp_elements(1014) <= cp_elements(1013);
    -- CP-element group 1015 fork  transition  place  input  bypass 
    -- predecessors 1014 
    -- successors 2310 2311 
    -- members (8) 
      -- 	branch_block_stmt_2042/if_stmt_3604_if_link/$exit
      -- 	branch_block_stmt_2042/if_stmt_3604_if_link/if_choice_transition
      -- 	branch_block_stmt_2042/iq_err_calcx_xexit_bb_58
      -- 	branch_block_stmt_2042/iq_err_calcx_xexit_bb_58_PhiReq/$entry
      -- 	branch_block_stmt_2042/iq_err_calcx_xexit_bb_58_PhiReq/phi_stmt_3626/$entry
      -- 	branch_block_stmt_2042/iq_err_calcx_xexit_bb_58_PhiReq/phi_stmt_3626/phi_stmt_3626_sources/$entry
      -- 	branch_block_stmt_2042/iq_err_calcx_xexit_bb_58_PhiReq/phi_stmt_3626/phi_stmt_3626_sources/type_cast_3629/$entry
      -- 	branch_block_stmt_2042/iq_err_calcx_xexit_bb_58_PhiReq/phi_stmt_3626/phi_stmt_3626_sources/type_cast_3629/SplitProtocol/$entry
      -- 
    if_choice_transition_14502_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_3604_branch_ack_1, ack => cp_elements(1015)); -- 
    -- CP-element group 1016 transition  bypass 
    -- predecessors 1013 
    -- successors 1017 
    -- members (1) 
      -- 	branch_block_stmt_2042/if_stmt_3604_else_link/$entry
      -- 
    cp_elements(1016) <= cp_elements(1013);
    -- CP-element group 1017 transition  place  input  bypass 
    -- predecessors 1016 
    -- successors 60 
    -- members (9) 
      -- 	branch_block_stmt_2042/if_stmt_3604_else_link/$exit
      -- 	branch_block_stmt_2042/if_stmt_3604_else_link/else_choice_transition
      -- 	branch_block_stmt_2042/iq_err_calcx_xexit_bb_56
      -- 	branch_block_stmt_2042/merge_stmt_3610_PhiReqMerge
      -- 	branch_block_stmt_2042/iq_err_calcx_xexit_bb_56_PhiReq/$entry
      -- 	branch_block_stmt_2042/iq_err_calcx_xexit_bb_56_PhiReq/$exit
      -- 	branch_block_stmt_2042/merge_stmt_3610_PhiAck/$entry
      -- 	branch_block_stmt_2042/merge_stmt_3610_PhiAck/$exit
      -- 	branch_block_stmt_2042/merge_stmt_3610_PhiAck/dummy
      -- 
    else_choice_transition_14506_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_3604_branch_ack_0, ack => cp_elements(1017)); -- 
    -- CP-element group 1018 fork  transition  bypass 
    -- predecessors 60 
    -- successors 1019 1020 
    -- members (1) 
      -- 	branch_block_stmt_2042/assign_stmt_3616/$entry
      -- 
    cp_elements(1018) <= cp_elements(60);
    -- CP-element group 1019 transition  output  bypass 
    -- predecessors 1018 
    -- successors 1022 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_3616/SGT_f32_u1_3615_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_3616/SGT_f32_u1_3615_Update/$entry
      -- 	branch_block_stmt_2042/assign_stmt_3616/SGT_f32_u1_3615_Update/cr
      -- 
    cp_elements(1019) <= cp_elements(1018);
    cr_14528_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1019), ack => SGT_f32_u1_3615_inst_req_1); -- 
    -- CP-element group 1020 transition  output  bypass 
    -- predecessors 1018 
    -- successors 1021 
    -- members (7) 
      -- 	branch_block_stmt_2042/assign_stmt_3616/SGT_f32_u1_3615_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_3616/R_iNsTr_85_3612_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_3616/R_iNsTr_85_3612_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3616/R_iNsTr_85_3612_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_3616/R_iNsTr_85_3612_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3616/SGT_f32_u1_3615_Sample/$entry
      -- 	branch_block_stmt_2042/assign_stmt_3616/SGT_f32_u1_3615_Sample/rr
      -- 
    cp_elements(1020) <= cp_elements(1018);
    rr_14523_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1020), ack => SGT_f32_u1_3615_inst_req_0); -- 
    -- CP-element group 1021 transition  input  bypass 
    -- predecessors 1020 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_3616/SGT_f32_u1_3615_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3616/SGT_f32_u1_3615_Sample/$exit
      -- 	branch_block_stmt_2042/assign_stmt_3616/SGT_f32_u1_3615_Sample/ra
      -- 
    ra_14524_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => SGT_f32_u1_3615_inst_ack_0, ack => cp_elements(1021)); -- 
    -- CP-element group 1022 branch  transition  place  input  bypass 
    -- predecessors 1019 
    -- successors 1023 1024 
    -- members (6) 
      -- 	branch_block_stmt_2042/if_stmt_3617__entry__
      -- 	branch_block_stmt_2042/assign_stmt_3616__exit__
      -- 	branch_block_stmt_2042/assign_stmt_3616/$exit
      -- 	branch_block_stmt_2042/assign_stmt_3616/SGT_f32_u1_3615_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3616/SGT_f32_u1_3615_Update/$exit
      -- 	branch_block_stmt_2042/assign_stmt_3616/SGT_f32_u1_3615_Update/ca
      -- 
    ca_14529_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => SGT_f32_u1_3615_inst_ack_1, ack => cp_elements(1022)); -- 
    -- CP-element group 1023 transition  place  dead  bypass 
    -- predecessors 1022 
    -- successors 61 
    -- members (8) 
      -- 	branch_block_stmt_2042/merge_stmt_3623__entry__
      -- 	branch_block_stmt_2042/if_stmt_3617__exit__
      -- 	branch_block_stmt_2042/if_stmt_3617_dead_link/$entry
      -- 	branch_block_stmt_2042/if_stmt_3617_dead_link/$exit
      -- 	branch_block_stmt_2042/if_stmt_3617_dead_link/dead_transition
      -- 	branch_block_stmt_2042/merge_stmt_3623_dead_link/$entry
      -- 	branch_block_stmt_2042/merge_stmt_3623_dead_link/$exit
      -- 	branch_block_stmt_2042/merge_stmt_3623_dead_link/dead_transition
      -- 
    cp_elements(1023) <= false;
    -- CP-element group 1024 transition  output  bypass 
    -- predecessors 1022 
    -- successors 1025 
    -- members (3) 
      -- 	branch_block_stmt_2042/if_stmt_3617_eval_test/$entry
      -- 	branch_block_stmt_2042/if_stmt_3617_eval_test/$exit
      -- 	branch_block_stmt_2042/if_stmt_3617_eval_test/branch_req
      -- 
    cp_elements(1024) <= cp_elements(1022);
    branch_req_14537_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1024), ack => if_stmt_3617_branch_req_0); -- 
    -- CP-element group 1025 branch  place  bypass 
    -- predecessors 1024 
    -- successors 1026 1028 
    -- members (1) 
      -- 	branch_block_stmt_2042/R_iNsTr_117_3618_place
      -- 
    cp_elements(1025) <= cp_elements(1024);
    -- CP-element group 1026 transition  bypass 
    -- predecessors 1025 
    -- successors 1027 
    -- members (1) 
      -- 	branch_block_stmt_2042/if_stmt_3617_if_link/$entry
      -- 
    cp_elements(1026) <= cp_elements(1025);
    -- CP-element group 1027 fork  transition  place  input  bypass 
    -- predecessors 1026 
    -- successors 2302 2303 
    -- members (8) 
      -- 	branch_block_stmt_2042/if_stmt_3617_if_link/$exit
      -- 	branch_block_stmt_2042/if_stmt_3617_if_link/if_choice_transition
      -- 	branch_block_stmt_2042/bb_56_bb_58
      -- 	branch_block_stmt_2042/bb_56_bb_58_PhiReq/$entry
      -- 	branch_block_stmt_2042/bb_56_bb_58_PhiReq/phi_stmt_3626/$entry
      -- 	branch_block_stmt_2042/bb_56_bb_58_PhiReq/phi_stmt_3626/phi_stmt_3626_sources/$entry
      -- 	branch_block_stmt_2042/bb_56_bb_58_PhiReq/phi_stmt_3626/phi_stmt_3626_sources/type_cast_3629/$entry
      -- 	branch_block_stmt_2042/bb_56_bb_58_PhiReq/phi_stmt_3626/phi_stmt_3626_sources/type_cast_3629/SplitProtocol/$entry
      -- 
    if_choice_transition_14542_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_3617_branch_ack_1, ack => cp_elements(1027)); -- 
    -- CP-element group 1028 transition  bypass 
    -- predecessors 1025 
    -- successors 1029 
    -- members (1) 
      -- 	branch_block_stmt_2042/if_stmt_3617_else_link/$entry
      -- 
    cp_elements(1028) <= cp_elements(1025);
    -- CP-element group 1029 transition  place  input  bypass 
    -- predecessors 1028 
    -- successors 61 
    -- members (9) 
      -- 	branch_block_stmt_2042/if_stmt_3617_else_link/$exit
      -- 	branch_block_stmt_2042/if_stmt_3617_else_link/else_choice_transition
      -- 	branch_block_stmt_2042/bb_56_bb_57
      -- 	branch_block_stmt_2042/merge_stmt_3623_PhiReqMerge
      -- 	branch_block_stmt_2042/bb_56_bb_57_PhiReq/$entry
      -- 	branch_block_stmt_2042/bb_56_bb_57_PhiReq/$exit
      -- 	branch_block_stmt_2042/merge_stmt_3623_PhiAck/$entry
      -- 	branch_block_stmt_2042/merge_stmt_3623_PhiAck/$exit
      -- 	branch_block_stmt_2042/merge_stmt_3623_PhiAck/dummy
      -- 
    else_choice_transition_14546_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_3617_branch_ack_0, ack => cp_elements(1029)); -- 
    -- CP-element group 1030 fork  transition  bypass 
    -- predecessors 2315 
    -- successors 1031 1032 1036 1037 1040 
    -- members (1) 
      -- 	branch_block_stmt_2042/assign_stmt_3642_to_assign_stmt_3653/$entry
      -- 
    cp_elements(1030) <= cp_elements(2315);
    -- CP-element group 1031 transition  output  bypass 
    -- predecessors 1030 
    -- successors 1034 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_3642_to_assign_stmt_3653/MUL_f32_f32_3641_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_3642_to_assign_stmt_3653/MUL_f32_f32_3641_Update/$entry
      -- 	branch_block_stmt_2042/assign_stmt_3642_to_assign_stmt_3653/MUL_f32_f32_3641_Update/cr
      -- 
    cp_elements(1031) <= cp_elements(1030);
    cr_14568_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1031), ack => MUL_f32_f32_3641_inst_req_1); -- 
    -- CP-element group 1032 transition  output  bypass 
    -- predecessors 1030 
    -- successors 1033 
    -- members (7) 
      -- 	branch_block_stmt_2042/assign_stmt_3642_to_assign_stmt_3653/MUL_f32_f32_3641_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_3642_to_assign_stmt_3653/R_iNsTr_82_3638_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_3642_to_assign_stmt_3653/R_iNsTr_82_3638_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3642_to_assign_stmt_3653/R_iNsTr_82_3638_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_3642_to_assign_stmt_3653/R_iNsTr_82_3638_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3642_to_assign_stmt_3653/MUL_f32_f32_3641_Sample/$entry
      -- 	branch_block_stmt_2042/assign_stmt_3642_to_assign_stmt_3653/MUL_f32_f32_3641_Sample/rr
      -- 
    cp_elements(1032) <= cp_elements(1030);
    rr_14563_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1032), ack => MUL_f32_f32_3641_inst_req_0); -- 
    -- CP-element group 1033 transition  input  bypass 
    -- predecessors 1032 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_3642_to_assign_stmt_3653/MUL_f32_f32_3641_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3642_to_assign_stmt_3653/MUL_f32_f32_3641_Sample/$exit
      -- 	branch_block_stmt_2042/assign_stmt_3642_to_assign_stmt_3653/MUL_f32_f32_3641_Sample/ra
      -- 
    ra_14564_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => MUL_f32_f32_3641_inst_ack_0, ack => cp_elements(1033)); -- 
    -- CP-element group 1034 transition  input  bypass 
    -- predecessors 1031 
    -- successors 1035 
    -- members (7) 
      -- 	branch_block_stmt_2042/assign_stmt_3642_to_assign_stmt_3653/MUL_f32_f32_3641_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3642_to_assign_stmt_3653/MUL_f32_f32_3641_Update/$exit
      -- 	branch_block_stmt_2042/assign_stmt_3642_to_assign_stmt_3653/MUL_f32_f32_3641_Update/ca
      -- 	branch_block_stmt_2042/assign_stmt_3642_to_assign_stmt_3653/R_iNsTr_113_3645_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_3642_to_assign_stmt_3653/R_iNsTr_113_3645_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3642_to_assign_stmt_3653/R_iNsTr_113_3645_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_3642_to_assign_stmt_3653/R_iNsTr_113_3645_update_completed_
      -- 
    ca_14569_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => MUL_f32_f32_3641_inst_ack_1, ack => cp_elements(1034)); -- 
    -- CP-element group 1035 join  transition  output  bypass 
    -- predecessors 1034 1037 
    -- successors 1038 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_3642_to_assign_stmt_3653/ADD_f32_f32_3646_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_3642_to_assign_stmt_3653/ADD_f32_f32_3646_Sample/$entry
      -- 	branch_block_stmt_2042/assign_stmt_3642_to_assign_stmt_3653/ADD_f32_f32_3646_Sample/rr
      -- 
    cp_element_group_1035: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1035"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1034) & cp_elements(1037);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1035), clk => clk, reset => reset); --
    end block;
    rr_14585_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1035), ack => ADD_f32_f32_3646_inst_req_0); -- 
    -- CP-element group 1036 transition  output  bypass 
    -- predecessors 1030 
    -- successors 1039 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_3642_to_assign_stmt_3653/ADD_f32_f32_3646_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_3642_to_assign_stmt_3653/ADD_f32_f32_3646_Update/$entry
      -- 	branch_block_stmt_2042/assign_stmt_3642_to_assign_stmt_3653/ADD_f32_f32_3646_Update/cr
      -- 
    cp_elements(1036) <= cp_elements(1030);
    cr_14590_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1036), ack => ADD_f32_f32_3646_inst_req_1); -- 
    -- CP-element group 1037 transition  bypass 
    -- predecessors 1030 
    -- successors 1035 
    -- members (4) 
      -- 	branch_block_stmt_2042/assign_stmt_3642_to_assign_stmt_3653/R_int_flux_errx_x1_3644_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_3642_to_assign_stmt_3653/R_int_flux_errx_x1_3644_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3642_to_assign_stmt_3653/R_int_flux_errx_x1_3644_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_3642_to_assign_stmt_3653/R_int_flux_errx_x1_3644_update_completed_
      -- 
    cp_elements(1037) <= cp_elements(1030);
    -- CP-element group 1038 transition  input  bypass 
    -- predecessors 1035 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_3642_to_assign_stmt_3653/ADD_f32_f32_3646_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3642_to_assign_stmt_3653/ADD_f32_f32_3646_Sample/$exit
      -- 	branch_block_stmt_2042/assign_stmt_3642_to_assign_stmt_3653/ADD_f32_f32_3646_Sample/ra
      -- 
    ra_14586_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_f32_f32_3646_inst_ack_0, ack => cp_elements(1038)); -- 
    -- CP-element group 1039 transition  input  output  bypass 
    -- predecessors 1036 
    -- successors 1041 
    -- members (10) 
      -- 	branch_block_stmt_2042/assign_stmt_3642_to_assign_stmt_3653/ADD_f32_f32_3646_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3642_to_assign_stmt_3653/ADD_f32_f32_3646_Update/$exit
      -- 	branch_block_stmt_2042/assign_stmt_3642_to_assign_stmt_3653/ADD_f32_f32_3646_Update/ca
      -- 	branch_block_stmt_2042/assign_stmt_3642_to_assign_stmt_3653/SLT_f32_u1_3652_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_3642_to_assign_stmt_3653/R_iNsTr_114_3649_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_3642_to_assign_stmt_3653/R_iNsTr_114_3649_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3642_to_assign_stmt_3653/R_iNsTr_114_3649_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_3642_to_assign_stmt_3653/R_iNsTr_114_3649_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3642_to_assign_stmt_3653/SLT_f32_u1_3652_Sample/$entry
      -- 	branch_block_stmt_2042/assign_stmt_3642_to_assign_stmt_3653/SLT_f32_u1_3652_Sample/rr
      -- 
    ca_14591_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_f32_f32_3646_inst_ack_1, ack => cp_elements(1039)); -- 
    rr_14603_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1039), ack => SLT_f32_u1_3652_inst_req_0); -- 
    -- CP-element group 1040 transition  output  bypass 
    -- predecessors 1030 
    -- successors 1042 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_3642_to_assign_stmt_3653/SLT_f32_u1_3652_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_3642_to_assign_stmt_3653/SLT_f32_u1_3652_Update/$entry
      -- 	branch_block_stmt_2042/assign_stmt_3642_to_assign_stmt_3653/SLT_f32_u1_3652_Update/cr
      -- 
    cp_elements(1040) <= cp_elements(1030);
    cr_14608_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1040), ack => SLT_f32_u1_3652_inst_req_1); -- 
    -- CP-element group 1041 transition  input  bypass 
    -- predecessors 1039 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_3642_to_assign_stmt_3653/SLT_f32_u1_3652_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3642_to_assign_stmt_3653/SLT_f32_u1_3652_Sample/$exit
      -- 	branch_block_stmt_2042/assign_stmt_3642_to_assign_stmt_3653/SLT_f32_u1_3652_Sample/ra
      -- 
    ra_14604_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => SLT_f32_u1_3652_inst_ack_0, ack => cp_elements(1041)); -- 
    -- CP-element group 1042 branch  transition  place  input  bypass 
    -- predecessors 1040 
    -- successors 1043 1044 
    -- members (6) 
      -- 	branch_block_stmt_2042/if_stmt_3654__entry__
      -- 	branch_block_stmt_2042/assign_stmt_3642_to_assign_stmt_3653__exit__
      -- 	branch_block_stmt_2042/assign_stmt_3642_to_assign_stmt_3653/$exit
      -- 	branch_block_stmt_2042/assign_stmt_3642_to_assign_stmt_3653/SLT_f32_u1_3652_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3642_to_assign_stmt_3653/SLT_f32_u1_3652_Update/$exit
      -- 	branch_block_stmt_2042/assign_stmt_3642_to_assign_stmt_3653/SLT_f32_u1_3652_Update/ca
      -- 
    ca_14609_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => SLT_f32_u1_3652_inst_ack_1, ack => cp_elements(1042)); -- 
    -- CP-element group 1043 transition  place  dead  bypass 
    -- predecessors 1042 
    -- successors 62 
    -- members (8) 
      -- 	branch_block_stmt_2042/merge_stmt_3660__entry__
      -- 	branch_block_stmt_2042/if_stmt_3654__exit__
      -- 	branch_block_stmt_2042/if_stmt_3654_dead_link/$entry
      -- 	branch_block_stmt_2042/if_stmt_3654_dead_link/$exit
      -- 	branch_block_stmt_2042/if_stmt_3654_dead_link/dead_transition
      -- 	branch_block_stmt_2042/merge_stmt_3660_dead_link/$entry
      -- 	branch_block_stmt_2042/merge_stmt_3660_dead_link/$exit
      -- 	branch_block_stmt_2042/merge_stmt_3660_dead_link/dead_transition
      -- 
    cp_elements(1043) <= false;
    -- CP-element group 1044 transition  output  bypass 
    -- predecessors 1042 
    -- successors 1045 
    -- members (3) 
      -- 	branch_block_stmt_2042/if_stmt_3654_eval_test/$entry
      -- 	branch_block_stmt_2042/if_stmt_3654_eval_test/$exit
      -- 	branch_block_stmt_2042/if_stmt_3654_eval_test/branch_req
      -- 
    cp_elements(1044) <= cp_elements(1042);
    branch_req_14617_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1044), ack => if_stmt_3654_branch_req_0); -- 
    -- CP-element group 1045 branch  place  bypass 
    -- predecessors 1044 
    -- successors 1046 1048 
    -- members (1) 
      -- 	branch_block_stmt_2042/R_iNsTr_115_3655_place
      -- 
    cp_elements(1045) <= cp_elements(1044);
    -- CP-element group 1046 transition  bypass 
    -- predecessors 1045 
    -- successors 1047 
    -- members (1) 
      -- 	branch_block_stmt_2042/if_stmt_3654_if_link/$entry
      -- 
    cp_elements(1046) <= cp_elements(1045);
    -- CP-element group 1047 fork  transition  place  input  bypass 
    -- predecessors 1046 
    -- successors 2316 2317 
    -- members (8) 
      -- 	branch_block_stmt_2042/if_stmt_3654_if_link/$exit
      -- 	branch_block_stmt_2042/if_stmt_3654_if_link/if_choice_transition
      -- 	branch_block_stmt_2042/bb_58_xx_xthread
      -- 	branch_block_stmt_2042/bb_58_xx_xthread_PhiReq/$entry
      -- 	branch_block_stmt_2042/bb_58_xx_xthread_PhiReq/phi_stmt_3687/$entry
      -- 	branch_block_stmt_2042/bb_58_xx_xthread_PhiReq/phi_stmt_3687/phi_stmt_3687_sources/$entry
      -- 	branch_block_stmt_2042/bb_58_xx_xthread_PhiReq/phi_stmt_3687/phi_stmt_3687_sources/type_cast_3690/$entry
      -- 	branch_block_stmt_2042/bb_58_xx_xthread_PhiReq/phi_stmt_3687/phi_stmt_3687_sources/type_cast_3690/SplitProtocol/$entry
      -- 
    if_choice_transition_14622_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_3654_branch_ack_1, ack => cp_elements(1047)); -- 
    -- CP-element group 1048 transition  bypass 
    -- predecessors 1045 
    -- successors 1049 
    -- members (1) 
      -- 	branch_block_stmt_2042/if_stmt_3654_else_link/$entry
      -- 
    cp_elements(1048) <= cp_elements(1045);
    -- CP-element group 1049 transition  place  input  bypass 
    -- predecessors 1048 
    -- successors 62 
    -- members (9) 
      -- 	branch_block_stmt_2042/if_stmt_3654_else_link/$exit
      -- 	branch_block_stmt_2042/if_stmt_3654_else_link/else_choice_transition
      -- 	branch_block_stmt_2042/bb_58_bb_59
      -- 	branch_block_stmt_2042/merge_stmt_3660_PhiReqMerge
      -- 	branch_block_stmt_2042/bb_58_bb_59_PhiReq/$entry
      -- 	branch_block_stmt_2042/bb_58_bb_59_PhiReq/$exit
      -- 	branch_block_stmt_2042/merge_stmt_3660_PhiAck/$entry
      -- 	branch_block_stmt_2042/merge_stmt_3660_PhiAck/$exit
      -- 	branch_block_stmt_2042/merge_stmt_3660_PhiAck/dummy
      -- 
    else_choice_transition_14626_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_3654_branch_ack_0, ack => cp_elements(1049)); -- 
    -- CP-element group 1050 fork  transition  bypass 
    -- predecessors 62 
    -- successors 1051 1052 
    -- members (1) 
      -- 	branch_block_stmt_2042/assign_stmt_3666/$entry
      -- 
    cp_elements(1050) <= cp_elements(62);
    -- CP-element group 1051 transition  output  bypass 
    -- predecessors 1050 
    -- successors 1054 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_3666/SGT_f32_u1_3665_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_3666/SGT_f32_u1_3665_Update/$entry
      -- 	branch_block_stmt_2042/assign_stmt_3666/SGT_f32_u1_3665_Update/cr
      -- 
    cp_elements(1051) <= cp_elements(1050);
    cr_14648_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1051), ack => SGT_f32_u1_3665_inst_req_1); -- 
    -- CP-element group 1052 transition  output  bypass 
    -- predecessors 1050 
    -- successors 1053 
    -- members (7) 
      -- 	branch_block_stmt_2042/assign_stmt_3666/SGT_f32_u1_3665_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_3666/R_iNsTr_114_3662_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_3666/R_iNsTr_114_3662_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3666/R_iNsTr_114_3662_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_3666/R_iNsTr_114_3662_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3666/SGT_f32_u1_3665_Sample/$entry
      -- 	branch_block_stmt_2042/assign_stmt_3666/SGT_f32_u1_3665_Sample/rr
      -- 
    cp_elements(1052) <= cp_elements(1050);
    rr_14643_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1052), ack => SGT_f32_u1_3665_inst_req_0); -- 
    -- CP-element group 1053 transition  input  bypass 
    -- predecessors 1052 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_3666/SGT_f32_u1_3665_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3666/SGT_f32_u1_3665_Sample/$exit
      -- 	branch_block_stmt_2042/assign_stmt_3666/SGT_f32_u1_3665_Sample/ra
      -- 
    ra_14644_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => SGT_f32_u1_3665_inst_ack_0, ack => cp_elements(1053)); -- 
    -- CP-element group 1054 branch  transition  place  input  bypass 
    -- predecessors 1051 
    -- successors 1055 1056 
    -- members (6) 
      -- 	branch_block_stmt_2042/if_stmt_3667__entry__
      -- 	branch_block_stmt_2042/assign_stmt_3666__exit__
      -- 	branch_block_stmt_2042/assign_stmt_3666/$exit
      -- 	branch_block_stmt_2042/assign_stmt_3666/SGT_f32_u1_3665_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3666/SGT_f32_u1_3665_Update/$exit
      -- 	branch_block_stmt_2042/assign_stmt_3666/SGT_f32_u1_3665_Update/ca
      -- 
    ca_14649_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => SGT_f32_u1_3665_inst_ack_1, ack => cp_elements(1054)); -- 
    -- CP-element group 1055 transition  place  dead  bypass 
    -- predecessors 1054 
    -- successors 63 
    -- members (8) 
      -- 	branch_block_stmt_2042/merge_stmt_3673__entry__
      -- 	branch_block_stmt_2042/if_stmt_3667__exit__
      -- 	branch_block_stmt_2042/if_stmt_3667_dead_link/$entry
      -- 	branch_block_stmt_2042/if_stmt_3667_dead_link/$exit
      -- 	branch_block_stmt_2042/if_stmt_3667_dead_link/dead_transition
      -- 	branch_block_stmt_2042/merge_stmt_3673_dead_link/$entry
      -- 	branch_block_stmt_2042/merge_stmt_3673_dead_link/$exit
      -- 	branch_block_stmt_2042/merge_stmt_3673_dead_link/dead_transition
      -- 
    cp_elements(1055) <= false;
    -- CP-element group 1056 transition  output  bypass 
    -- predecessors 1054 
    -- successors 1057 
    -- members (3) 
      -- 	branch_block_stmt_2042/if_stmt_3667_eval_test/$entry
      -- 	branch_block_stmt_2042/if_stmt_3667_eval_test/$exit
      -- 	branch_block_stmt_2042/if_stmt_3667_eval_test/branch_req
      -- 
    cp_elements(1056) <= cp_elements(1054);
    branch_req_14657_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1056), ack => if_stmt_3667_branch_req_0); -- 
    -- CP-element group 1057 branch  place  bypass 
    -- predecessors 1056 
    -- successors 1058 1060 
    -- members (1) 
      -- 	branch_block_stmt_2042/R_iNsTr_151_3668_place
      -- 
    cp_elements(1057) <= cp_elements(1056);
    -- CP-element group 1058 transition  bypass 
    -- predecessors 1057 
    -- successors 1059 
    -- members (1) 
      -- 	branch_block_stmt_2042/if_stmt_3667_if_link/$entry
      -- 
    cp_elements(1058) <= cp_elements(1057);
    -- CP-element group 1059 fork  transition  place  input  bypass 
    -- predecessors 1058 
    -- successors 2319 2320 
    -- members (8) 
      -- 	branch_block_stmt_2042/if_stmt_3667_if_link/$exit
      -- 	branch_block_stmt_2042/if_stmt_3667_if_link/if_choice_transition
      -- 	branch_block_stmt_2042/bb_59_xx_xthread
      -- 	branch_block_stmt_2042/bb_59_xx_xthread_PhiReq/$entry
      -- 	branch_block_stmt_2042/bb_59_xx_xthread_PhiReq/phi_stmt_3687/$entry
      -- 	branch_block_stmt_2042/bb_59_xx_xthread_PhiReq/phi_stmt_3687/phi_stmt_3687_sources/$entry
      -- 	branch_block_stmt_2042/bb_59_xx_xthread_PhiReq/phi_stmt_3687/phi_stmt_3687_sources/type_cast_3690/$entry
      -- 	branch_block_stmt_2042/bb_59_xx_xthread_PhiReq/phi_stmt_3687/phi_stmt_3687_sources/type_cast_3690/SplitProtocol/$entry
      -- 
    if_choice_transition_14662_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_3667_branch_ack_1, ack => cp_elements(1059)); -- 
    -- CP-element group 1060 transition  bypass 
    -- predecessors 1057 
    -- successors 1061 
    -- members (1) 
      -- 	branch_block_stmt_2042/if_stmt_3667_else_link/$entry
      -- 
    cp_elements(1060) <= cp_elements(1057);
    -- CP-element group 1061 transition  place  input  bypass 
    -- predecessors 1060 
    -- successors 63 
    -- members (9) 
      -- 	branch_block_stmt_2042/if_stmt_3667_else_link/$exit
      -- 	branch_block_stmt_2042/if_stmt_3667_else_link/else_choice_transition
      -- 	branch_block_stmt_2042/bb_59_bb_60
      -- 	branch_block_stmt_2042/merge_stmt_3673_PhiReqMerge
      -- 	branch_block_stmt_2042/bb_59_bb_60_PhiReq/$entry
      -- 	branch_block_stmt_2042/bb_59_bb_60_PhiReq/$exit
      -- 	branch_block_stmt_2042/merge_stmt_3673_PhiAck/$entry
      -- 	branch_block_stmt_2042/merge_stmt_3673_PhiAck/$exit
      -- 	branch_block_stmt_2042/merge_stmt_3673_PhiAck/dummy
      -- 
    else_choice_transition_14666_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_3667_branch_ack_0, ack => cp_elements(1061)); -- 
    -- CP-element group 1062 fork  transition  bypass 
    -- predecessors 63 
    -- successors 1063 1064 
    -- members (1) 
      -- 	branch_block_stmt_2042/assign_stmt_3679/$entry
      -- 
    cp_elements(1062) <= cp_elements(63);
    -- CP-element group 1063 transition  output  bypass 
    -- predecessors 1062 
    -- successors 1066 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_3679/EQ_f32_u1_3678_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_3679/EQ_f32_u1_3678_Update/$entry
      -- 	branch_block_stmt_2042/assign_stmt_3679/EQ_f32_u1_3678_Update/cr
      -- 
    cp_elements(1063) <= cp_elements(1062);
    cr_14688_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1063), ack => EQ_f32_u1_3678_inst_req_1); -- 
    -- CP-element group 1064 transition  output  bypass 
    -- predecessors 1062 
    -- successors 1065 
    -- members (7) 
      -- 	branch_block_stmt_2042/assign_stmt_3679/EQ_f32_u1_3678_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_3679/R_iNsTr_114_3675_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_3679/R_iNsTr_114_3675_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3679/R_iNsTr_114_3675_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_3679/R_iNsTr_114_3675_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3679/EQ_f32_u1_3678_Sample/$entry
      -- 	branch_block_stmt_2042/assign_stmt_3679/EQ_f32_u1_3678_Sample/rr
      -- 
    cp_elements(1064) <= cp_elements(1062);
    rr_14683_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1064), ack => EQ_f32_u1_3678_inst_req_0); -- 
    -- CP-element group 1065 transition  input  bypass 
    -- predecessors 1064 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_3679/EQ_f32_u1_3678_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3679/EQ_f32_u1_3678_Sample/$exit
      -- 	branch_block_stmt_2042/assign_stmt_3679/EQ_f32_u1_3678_Sample/ra
      -- 
    ra_14684_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_f32_u1_3678_inst_ack_0, ack => cp_elements(1065)); -- 
    -- CP-element group 1066 branch  transition  place  input  bypass 
    -- predecessors 1063 
    -- successors 1067 1068 
    -- members (6) 
      -- 	branch_block_stmt_2042/assign_stmt_3679__exit__
      -- 	branch_block_stmt_2042/if_stmt_3680__entry__
      -- 	branch_block_stmt_2042/assign_stmt_3679/$exit
      -- 	branch_block_stmt_2042/assign_stmt_3679/EQ_f32_u1_3678_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3679/EQ_f32_u1_3678_Update/$exit
      -- 	branch_block_stmt_2042/assign_stmt_3679/EQ_f32_u1_3678_Update/ca
      -- 
    ca_14689_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_f32_u1_3678_inst_ack_1, ack => cp_elements(1066)); -- 
    -- CP-element group 1067 transition  place  dead  bypass 
    -- predecessors 1066 
    -- successors 64 
    -- members (8) 
      -- 	branch_block_stmt_2042/merge_stmt_3686__entry__
      -- 	branch_block_stmt_2042/if_stmt_3680__exit__
      -- 	branch_block_stmt_2042/if_stmt_3680_dead_link/$entry
      -- 	branch_block_stmt_2042/if_stmt_3680_dead_link/$exit
      -- 	branch_block_stmt_2042/if_stmt_3680_dead_link/dead_transition
      -- 	branch_block_stmt_2042/merge_stmt_3686_dead_link/$entry
      -- 	branch_block_stmt_2042/merge_stmt_3686_dead_link/$exit
      -- 	branch_block_stmt_2042/merge_stmt_3686_dead_link/dead_transition
      -- 
    cp_elements(1067) <= false;
    -- CP-element group 1068 transition  output  bypass 
    -- predecessors 1066 
    -- successors 1069 
    -- members (3) 
      -- 	branch_block_stmt_2042/if_stmt_3680_eval_test/$entry
      -- 	branch_block_stmt_2042/if_stmt_3680_eval_test/$exit
      -- 	branch_block_stmt_2042/if_stmt_3680_eval_test/branch_req
      -- 
    cp_elements(1068) <= cp_elements(1066);
    branch_req_14697_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1068), ack => if_stmt_3680_branch_req_0); -- 
    -- CP-element group 1069 branch  place  bypass 
    -- predecessors 1068 
    -- successors 1070 1072 
    -- members (1) 
      -- 	branch_block_stmt_2042/R_iNsTr_186_3681_place
      -- 
    cp_elements(1069) <= cp_elements(1068);
    -- CP-element group 1070 transition  bypass 
    -- predecessors 1069 
    -- successors 1071 
    -- members (1) 
      -- 	branch_block_stmt_2042/if_stmt_3680_if_link/$entry
      -- 
    cp_elements(1070) <= cp_elements(1069);
    -- CP-element group 1071 fork  transition  place  input  bypass 
    -- predecessors 1070 
    -- successors 2575 2576 
    -- members (8) 
      -- 	branch_block_stmt_2042/if_stmt_3680_if_link/$exit
      -- 	branch_block_stmt_2042/if_stmt_3680_if_link/if_choice_transition
      -- 	branch_block_stmt_2042/bb_60_fdiv32x_xexit
      -- 	branch_block_stmt_2042/bb_60_fdiv32x_xexit_PhiReq/$entry
      -- 	branch_block_stmt_2042/bb_60_fdiv32x_xexit_PhiReq/phi_stmt_4035/$entry
      -- 	branch_block_stmt_2042/bb_60_fdiv32x_xexit_PhiReq/phi_stmt_4035/phi_stmt_4035_sources/$entry
      -- 	branch_block_stmt_2042/bb_60_fdiv32x_xexit_PhiReq/phi_stmt_4035/phi_stmt_4035_sources/type_cast_4038/$entry
      -- 	branch_block_stmt_2042/bb_60_fdiv32x_xexit_PhiReq/phi_stmt_4035/phi_stmt_4035_sources/type_cast_4038/SplitProtocol/$entry
      -- 
    if_choice_transition_14702_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_3680_branch_ack_1, ack => cp_elements(1071)); -- 
    -- CP-element group 1072 transition  bypass 
    -- predecessors 1069 
    -- successors 1073 
    -- members (1) 
      -- 	branch_block_stmt_2042/if_stmt_3680_else_link/$entry
      -- 
    cp_elements(1072) <= cp_elements(1069);
    -- CP-element group 1073 fork  transition  place  input  bypass 
    -- predecessors 1072 
    -- successors 2322 2324 
    -- members (8) 
      -- 	branch_block_stmt_2042/if_stmt_3680_else_link/$exit
      -- 	branch_block_stmt_2042/if_stmt_3680_else_link/else_choice_transition
      -- 	branch_block_stmt_2042/bb_60_xx_xthread
      -- 	branch_block_stmt_2042/bb_60_xx_xthread_PhiReq/$entry
      -- 	branch_block_stmt_2042/bb_60_xx_xthread_PhiReq/phi_stmt_3687/$entry
      -- 	branch_block_stmt_2042/bb_60_xx_xthread_PhiReq/phi_stmt_3687/phi_stmt_3687_sources/$entry
      -- 	branch_block_stmt_2042/bb_60_xx_xthread_PhiReq/phi_stmt_3687/phi_stmt_3687_sources/type_cast_3690/$entry
      -- 	branch_block_stmt_2042/bb_60_xx_xthread_PhiReq/phi_stmt_3687/phi_stmt_3687_sources/type_cast_3690/SplitProtocol/$entry
      -- 
    else_choice_transition_14706_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_3680_branch_ack_0, ack => cp_elements(1073)); -- 
    -- CP-element group 1074 fork  transition  bypass 
    -- predecessors 64 
    -- successors 1075 1076 1079 1082 1085 
    -- members (1) 
      -- 	branch_block_stmt_2042/assign_stmt_3701_to_assign_stmt_3719/$entry
      -- 
    cp_elements(1074) <= cp_elements(64);
    -- CP-element group 1075 transition  output  bypass 
    -- predecessors 1074 
    -- successors 1078 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_3701_to_assign_stmt_3719/type_cast_3700_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_3701_to_assign_stmt_3719/type_cast_3700_Update/$entry
      -- 	branch_block_stmt_2042/assign_stmt_3701_to_assign_stmt_3719/type_cast_3700_Update/cr
      -- 
    cp_elements(1075) <= cp_elements(1074);
    cr_14728_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1075), ack => type_cast_3700_inst_req_1); -- 
    -- CP-element group 1076 transition  output  bypass 
    -- predecessors 1074 
    -- successors 1077 
    -- members (7) 
      -- 	branch_block_stmt_2042/assign_stmt_3701_to_assign_stmt_3719/type_cast_3700_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_3701_to_assign_stmt_3719/R_tmp10x_xi55x_xin_3699_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_3701_to_assign_stmt_3719/R_tmp10x_xi55x_xin_3699_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3701_to_assign_stmt_3719/R_tmp10x_xi55x_xin_3699_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_3701_to_assign_stmt_3719/R_tmp10x_xi55x_xin_3699_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3701_to_assign_stmt_3719/type_cast_3700_Sample/$entry
      -- 	branch_block_stmt_2042/assign_stmt_3701_to_assign_stmt_3719/type_cast_3700_Sample/rr
      -- 
    cp_elements(1076) <= cp_elements(1074);
    rr_14723_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1076), ack => type_cast_3700_inst_req_0); -- 
    -- CP-element group 1077 transition  input  bypass 
    -- predecessors 1076 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_3701_to_assign_stmt_3719/type_cast_3700_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3701_to_assign_stmt_3719/type_cast_3700_Sample/$exit
      -- 	branch_block_stmt_2042/assign_stmt_3701_to_assign_stmt_3719/type_cast_3700_Sample/ra
      -- 
    ra_14724_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3700_inst_ack_0, ack => cp_elements(1077)); -- 
    -- CP-element group 1078 transition  input  output  bypass 
    -- predecessors 1075 
    -- successors 1080 
    -- members (10) 
      -- 	branch_block_stmt_2042/assign_stmt_3701_to_assign_stmt_3719/type_cast_3700_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3701_to_assign_stmt_3719/type_cast_3700_Update/$exit
      -- 	branch_block_stmt_2042/assign_stmt_3701_to_assign_stmt_3719/type_cast_3700_Update/ca
      -- 	branch_block_stmt_2042/assign_stmt_3701_to_assign_stmt_3719/SHL_u32_u32_3706_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_3701_to_assign_stmt_3719/R_tmp10x_xi55_3703_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_3701_to_assign_stmt_3719/R_tmp10x_xi55_3703_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3701_to_assign_stmt_3719/R_tmp10x_xi55_3703_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_3701_to_assign_stmt_3719/R_tmp10x_xi55_3703_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3701_to_assign_stmt_3719/SHL_u32_u32_3706_Sample/$entry
      -- 	branch_block_stmt_2042/assign_stmt_3701_to_assign_stmt_3719/SHL_u32_u32_3706_Sample/rr
      -- 
    ca_14729_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3700_inst_ack_1, ack => cp_elements(1078)); -- 
    rr_14741_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1078), ack => SHL_u32_u32_3706_inst_req_0); -- 
    -- CP-element group 1079 transition  output  bypass 
    -- predecessors 1074 
    -- successors 1081 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_3701_to_assign_stmt_3719/SHL_u32_u32_3706_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_3701_to_assign_stmt_3719/SHL_u32_u32_3706_Update/$entry
      -- 	branch_block_stmt_2042/assign_stmt_3701_to_assign_stmt_3719/SHL_u32_u32_3706_Update/cr
      -- 
    cp_elements(1079) <= cp_elements(1074);
    cr_14746_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1079), ack => SHL_u32_u32_3706_inst_req_1); -- 
    -- CP-element group 1080 transition  input  bypass 
    -- predecessors 1078 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_3701_to_assign_stmt_3719/SHL_u32_u32_3706_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3701_to_assign_stmt_3719/SHL_u32_u32_3706_Sample/$exit
      -- 	branch_block_stmt_2042/assign_stmt_3701_to_assign_stmt_3719/SHL_u32_u32_3706_Sample/ra
      -- 
    ra_14742_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => SHL_u32_u32_3706_inst_ack_0, ack => cp_elements(1080)); -- 
    -- CP-element group 1081 transition  input  output  bypass 
    -- predecessors 1079 
    -- successors 1083 
    -- members (10) 
      -- 	branch_block_stmt_2042/assign_stmt_3701_to_assign_stmt_3719/SHL_u32_u32_3706_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3701_to_assign_stmt_3719/SHL_u32_u32_3706_Update/$exit
      -- 	branch_block_stmt_2042/assign_stmt_3701_to_assign_stmt_3719/SHL_u32_u32_3706_Update/ca
      -- 	branch_block_stmt_2042/assign_stmt_3701_to_assign_stmt_3719/AND_u32_u32_3712_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_3701_to_assign_stmt_3719/R_iNsTr_147_3709_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_3701_to_assign_stmt_3719/R_iNsTr_147_3709_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3701_to_assign_stmt_3719/R_iNsTr_147_3709_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_3701_to_assign_stmt_3719/R_iNsTr_147_3709_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3701_to_assign_stmt_3719/AND_u32_u32_3712_Sample/$entry
      -- 	branch_block_stmt_2042/assign_stmt_3701_to_assign_stmt_3719/AND_u32_u32_3712_Sample/rr
      -- 
    ca_14747_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => SHL_u32_u32_3706_inst_ack_1, ack => cp_elements(1081)); -- 
    rr_14759_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1081), ack => AND_u32_u32_3712_inst_req_0); -- 
    -- CP-element group 1082 transition  output  bypass 
    -- predecessors 1074 
    -- successors 1084 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_3701_to_assign_stmt_3719/AND_u32_u32_3712_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_3701_to_assign_stmt_3719/AND_u32_u32_3712_Update/$entry
      -- 	branch_block_stmt_2042/assign_stmt_3701_to_assign_stmt_3719/AND_u32_u32_3712_Update/cr
      -- 
    cp_elements(1082) <= cp_elements(1074);
    cr_14764_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1082), ack => AND_u32_u32_3712_inst_req_1); -- 
    -- CP-element group 1083 transition  input  bypass 
    -- predecessors 1081 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_3701_to_assign_stmt_3719/AND_u32_u32_3712_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3701_to_assign_stmt_3719/AND_u32_u32_3712_Sample/$exit
      -- 	branch_block_stmt_2042/assign_stmt_3701_to_assign_stmt_3719/AND_u32_u32_3712_Sample/ra
      -- 
    ra_14760_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => AND_u32_u32_3712_inst_ack_0, ack => cp_elements(1083)); -- 
    -- CP-element group 1084 transition  input  output  bypass 
    -- predecessors 1082 
    -- successors 1086 
    -- members (10) 
      -- 	branch_block_stmt_2042/assign_stmt_3701_to_assign_stmt_3719/AND_u32_u32_3712_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3701_to_assign_stmt_3719/AND_u32_u32_3712_Update/$exit
      -- 	branch_block_stmt_2042/assign_stmt_3701_to_assign_stmt_3719/AND_u32_u32_3712_Update/ca
      -- 	branch_block_stmt_2042/assign_stmt_3701_to_assign_stmt_3719/OR_u32_u32_3718_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_3701_to_assign_stmt_3719/R_iNsTr_148_3715_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_3701_to_assign_stmt_3719/R_iNsTr_148_3715_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3701_to_assign_stmt_3719/R_iNsTr_148_3715_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_3701_to_assign_stmt_3719/R_iNsTr_148_3715_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3701_to_assign_stmt_3719/OR_u32_u32_3718_Sample/$entry
      -- 	branch_block_stmt_2042/assign_stmt_3701_to_assign_stmt_3719/OR_u32_u32_3718_Sample/rr
      -- 
    ca_14765_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => AND_u32_u32_3712_inst_ack_1, ack => cp_elements(1084)); -- 
    rr_14777_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1084), ack => OR_u32_u32_3718_inst_req_0); -- 
    -- CP-element group 1085 transition  output  bypass 
    -- predecessors 1074 
    -- successors 1087 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_3701_to_assign_stmt_3719/OR_u32_u32_3718_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_3701_to_assign_stmt_3719/OR_u32_u32_3718_Update/$entry
      -- 	branch_block_stmt_2042/assign_stmt_3701_to_assign_stmt_3719/OR_u32_u32_3718_Update/cr
      -- 
    cp_elements(1085) <= cp_elements(1074);
    cr_14782_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1085), ack => OR_u32_u32_3718_inst_req_1); -- 
    -- CP-element group 1086 transition  input  bypass 
    -- predecessors 1084 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_3701_to_assign_stmt_3719/OR_u32_u32_3718_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3701_to_assign_stmt_3719/OR_u32_u32_3718_Sample/$exit
      -- 	branch_block_stmt_2042/assign_stmt_3701_to_assign_stmt_3719/OR_u32_u32_3718_Sample/ra
      -- 
    ra_14778_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => OR_u32_u32_3718_inst_ack_0, ack => cp_elements(1086)); -- 
    -- CP-element group 1087 transition  place  input  bypass 
    -- predecessors 1085 
    -- successors 2350 
    -- members (6) 
      -- 	branch_block_stmt_2042/assign_stmt_3701_to_assign_stmt_3719__exit__
      -- 	branch_block_stmt_2042/xx_xthread_bbx_xnph7x_xix_xi
      -- 	branch_block_stmt_2042/assign_stmt_3701_to_assign_stmt_3719/$exit
      -- 	branch_block_stmt_2042/assign_stmt_3701_to_assign_stmt_3719/OR_u32_u32_3718_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3701_to_assign_stmt_3719/OR_u32_u32_3718_Update/$exit
      -- 	branch_block_stmt_2042/assign_stmt_3701_to_assign_stmt_3719/OR_u32_u32_3718_Update/ca
      -- 
    ca_14783_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => OR_u32_u32_3718_inst_ack_1, ack => cp_elements(1087)); -- 
    -- CP-element group 1088 fork  transition  bypass 
    -- predecessors 65 
    -- successors 1089 1090 1093 
    -- members (1) 
      -- 	branch_block_stmt_2042/assign_stmt_3741_to_assign_stmt_3747/$entry
      -- 
    cp_elements(1088) <= cp_elements(65);
    -- CP-element group 1089 transition  output  bypass 
    -- predecessors 1088 
    -- successors 1092 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_3741_to_assign_stmt_3747/LSHR_u32_u32_3740_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_3741_to_assign_stmt_3747/LSHR_u32_u32_3740_Update/$entry
      -- 	branch_block_stmt_2042/assign_stmt_3741_to_assign_stmt_3747/LSHR_u32_u32_3740_Update/cr
      -- 
    cp_elements(1089) <= cp_elements(1088);
    cr_14803_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1089), ack => LSHR_u32_u32_3740_inst_req_1); -- 
    -- CP-element group 1090 transition  output  bypass 
    -- predecessors 1088 
    -- successors 1091 
    -- members (7) 
      -- 	branch_block_stmt_2042/assign_stmt_3741_to_assign_stmt_3747/LSHR_u32_u32_3740_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_3741_to_assign_stmt_3747/R_xx_x016x_xix_xi_3737_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_3741_to_assign_stmt_3747/R_xx_x016x_xix_xi_3737_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3741_to_assign_stmt_3747/R_xx_x016x_xix_xi_3737_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_3741_to_assign_stmt_3747/R_xx_x016x_xix_xi_3737_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3741_to_assign_stmt_3747/LSHR_u32_u32_3740_Sample/$entry
      -- 	branch_block_stmt_2042/assign_stmt_3741_to_assign_stmt_3747/LSHR_u32_u32_3740_Sample/rr
      -- 
    cp_elements(1090) <= cp_elements(1088);
    rr_14798_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1090), ack => LSHR_u32_u32_3740_inst_req_0); -- 
    -- CP-element group 1091 transition  input  bypass 
    -- predecessors 1090 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_3741_to_assign_stmt_3747/LSHR_u32_u32_3740_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3741_to_assign_stmt_3747/LSHR_u32_u32_3740_Sample/$exit
      -- 	branch_block_stmt_2042/assign_stmt_3741_to_assign_stmt_3747/LSHR_u32_u32_3740_Sample/ra
      -- 
    ra_14799_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => LSHR_u32_u32_3740_inst_ack_0, ack => cp_elements(1091)); -- 
    -- CP-element group 1092 transition  input  output  bypass 
    -- predecessors 1089 
    -- successors 1094 
    -- members (10) 
      -- 	branch_block_stmt_2042/assign_stmt_3741_to_assign_stmt_3747/LSHR_u32_u32_3740_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3741_to_assign_stmt_3747/LSHR_u32_u32_3740_Update/$exit
      -- 	branch_block_stmt_2042/assign_stmt_3741_to_assign_stmt_3747/LSHR_u32_u32_3740_Update/ca
      -- 	branch_block_stmt_2042/assign_stmt_3741_to_assign_stmt_3747/UGT_u32_u1_3746_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_3741_to_assign_stmt_3747/R_iNsTr_183_3743_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_3741_to_assign_stmt_3747/R_iNsTr_183_3743_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3741_to_assign_stmt_3747/R_iNsTr_183_3743_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_3741_to_assign_stmt_3747/R_iNsTr_183_3743_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3741_to_assign_stmt_3747/UGT_u32_u1_3746_Sample/$entry
      -- 	branch_block_stmt_2042/assign_stmt_3741_to_assign_stmt_3747/UGT_u32_u1_3746_Sample/rr
      -- 
    ca_14804_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => LSHR_u32_u32_3740_inst_ack_1, ack => cp_elements(1092)); -- 
    rr_14816_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1092), ack => UGT_u32_u1_3746_inst_req_0); -- 
    -- CP-element group 1093 transition  output  bypass 
    -- predecessors 1088 
    -- successors 1095 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_3741_to_assign_stmt_3747/UGT_u32_u1_3746_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_3741_to_assign_stmt_3747/UGT_u32_u1_3746_Update/$entry
      -- 	branch_block_stmt_2042/assign_stmt_3741_to_assign_stmt_3747/UGT_u32_u1_3746_Update/cr
      -- 
    cp_elements(1093) <= cp_elements(1088);
    cr_14821_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1093), ack => UGT_u32_u1_3746_inst_req_1); -- 
    -- CP-element group 1094 transition  input  bypass 
    -- predecessors 1092 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_3741_to_assign_stmt_3747/UGT_u32_u1_3746_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3741_to_assign_stmt_3747/UGT_u32_u1_3746_Sample/$exit
      -- 	branch_block_stmt_2042/assign_stmt_3741_to_assign_stmt_3747/UGT_u32_u1_3746_Sample/ra
      -- 
    ra_14817_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => UGT_u32_u1_3746_inst_ack_0, ack => cp_elements(1094)); -- 
    -- CP-element group 1095 branch  transition  place  input  bypass 
    -- predecessors 1093 
    -- successors 1096 1097 
    -- members (6) 
      -- 	branch_block_stmt_2042/assign_stmt_3741_to_assign_stmt_3747__exit__
      -- 	branch_block_stmt_2042/if_stmt_3748__entry__
      -- 	branch_block_stmt_2042/assign_stmt_3741_to_assign_stmt_3747/$exit
      -- 	branch_block_stmt_2042/assign_stmt_3741_to_assign_stmt_3747/UGT_u32_u1_3746_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3741_to_assign_stmt_3747/UGT_u32_u1_3746_Update/$exit
      -- 	branch_block_stmt_2042/assign_stmt_3741_to_assign_stmt_3747/UGT_u32_u1_3746_Update/ca
      -- 
    ca_14822_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => UGT_u32_u1_3746_inst_ack_1, ack => cp_elements(1095)); -- 
    -- CP-element group 1096 transition  place  dead  bypass 
    -- predecessors 1095 
    -- successors 66 
    -- members (8) 
      -- 	branch_block_stmt_2042/if_stmt_3748__exit__
      -- 	branch_block_stmt_2042/merge_stmt_3754__entry__
      -- 	branch_block_stmt_2042/if_stmt_3748_dead_link/$entry
      -- 	branch_block_stmt_2042/if_stmt_3748_dead_link/$exit
      -- 	branch_block_stmt_2042/if_stmt_3748_dead_link/dead_transition
      -- 	branch_block_stmt_2042/merge_stmt_3754_dead_link/$entry
      -- 	branch_block_stmt_2042/merge_stmt_3754_dead_link/$exit
      -- 	branch_block_stmt_2042/merge_stmt_3754_dead_link/dead_transition
      -- 
    cp_elements(1096) <= false;
    -- CP-element group 1097 transition  output  bypass 
    -- predecessors 1095 
    -- successors 1098 
    -- members (3) 
      -- 	branch_block_stmt_2042/if_stmt_3748_eval_test/$entry
      -- 	branch_block_stmt_2042/if_stmt_3748_eval_test/$exit
      -- 	branch_block_stmt_2042/if_stmt_3748_eval_test/branch_req
      -- 
    cp_elements(1097) <= cp_elements(1095);
    branch_req_14830_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1097), ack => if_stmt_3748_branch_req_0); -- 
    -- CP-element group 1098 branch  place  bypass 
    -- predecessors 1097 
    -- successors 1099 1101 
    -- members (1) 
      -- 	branch_block_stmt_2042/R_iNsTr_184_3749_place
      -- 
    cp_elements(1098) <= cp_elements(1097);
    -- CP-element group 1099 transition  bypass 
    -- predecessors 1098 
    -- successors 1100 
    -- members (1) 
      -- 	branch_block_stmt_2042/if_stmt_3748_if_link/$entry
      -- 
    cp_elements(1099) <= cp_elements(1098);
    -- CP-element group 1100 transition  place  input  bypass 
    -- predecessors 1099 
    -- successors 66 
    -- members (9) 
      -- 	branch_block_stmt_2042/if_stmt_3748_if_link/$exit
      -- 	branch_block_stmt_2042/if_stmt_3748_if_link/if_choice_transition
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xi_bbx_xnphx_xix_xix_xpreheader
      -- 	branch_block_stmt_2042/merge_stmt_3754_PhiReqMerge
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xi_bbx_xnphx_xix_xix_xpreheader_PhiReq/$entry
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xi_bbx_xnphx_xix_xix_xpreheader_PhiReq/$exit
      -- 	branch_block_stmt_2042/merge_stmt_3754_PhiAck/$entry
      -- 	branch_block_stmt_2042/merge_stmt_3754_PhiAck/$exit
      -- 	branch_block_stmt_2042/merge_stmt_3754_PhiAck/dummy
      -- 
    if_choice_transition_14835_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_3748_branch_ack_1, ack => cp_elements(1100)); -- 
    -- CP-element group 1101 transition  bypass 
    -- predecessors 1098 
    -- successors 1102 
    -- members (1) 
      -- 	branch_block_stmt_2042/if_stmt_3748_else_link/$entry
      -- 
    cp_elements(1101) <= cp_elements(1098);
    -- CP-element group 1102 transition  place  input  bypass 
    -- predecessors 1101 
    -- successors 2421 
    -- members (3) 
      -- 	branch_block_stmt_2042/if_stmt_3748_else_link/$exit
      -- 	branch_block_stmt_2042/if_stmt_3748_else_link/else_choice_transition
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xi_xx_x_crit_edgex_xix_xi
      -- 
    else_choice_transition_14839_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_3748_branch_ack_0, ack => cp_elements(1102)); -- 
    -- CP-element group 1103 fork  transition  bypass 
    -- predecessors 67 
    -- successors 1104 1105 1108 1109 1113 1114 
    -- members (1) 
      -- 	branch_block_stmt_2042/assign_stmt_3777_to_assign_stmt_3788/$entry
      -- 
    cp_elements(1103) <= cp_elements(67);
    -- CP-element group 1104 transition  output  bypass 
    -- predecessors 1103 
    -- successors 1107 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_3777_to_assign_stmt_3788/SHL_u32_u32_3776_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_3777_to_assign_stmt_3788/SHL_u32_u32_3776_Update/$entry
      -- 	branch_block_stmt_2042/assign_stmt_3777_to_assign_stmt_3788/SHL_u32_u32_3776_Update/cr
      -- 
    cp_elements(1104) <= cp_elements(1103);
    cr_14861_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1104), ack => SHL_u32_u32_3776_inst_req_1); -- 
    -- CP-element group 1105 transition  output  bypass 
    -- predecessors 1103 
    -- successors 1106 
    -- members (7) 
      -- 	branch_block_stmt_2042/assign_stmt_3777_to_assign_stmt_3788/SHL_u32_u32_3776_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_3777_to_assign_stmt_3788/R_shifted_divisorx_x03x_xix_xi_3773_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_3777_to_assign_stmt_3788/R_shifted_divisorx_x03x_xix_xi_3773_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3777_to_assign_stmt_3788/R_shifted_divisorx_x03x_xix_xi_3773_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_3777_to_assign_stmt_3788/R_shifted_divisorx_x03x_xix_xi_3773_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3777_to_assign_stmt_3788/SHL_u32_u32_3776_Sample/$entry
      -- 	branch_block_stmt_2042/assign_stmt_3777_to_assign_stmt_3788/SHL_u32_u32_3776_Sample/rr
      -- 
    cp_elements(1105) <= cp_elements(1103);
    rr_14856_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1105), ack => SHL_u32_u32_3776_inst_req_0); -- 
    -- CP-element group 1106 transition  input  bypass 
    -- predecessors 1105 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_3777_to_assign_stmt_3788/SHL_u32_u32_3776_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3777_to_assign_stmt_3788/SHL_u32_u32_3776_Sample/$exit
      -- 	branch_block_stmt_2042/assign_stmt_3777_to_assign_stmt_3788/SHL_u32_u32_3776_Sample/ra
      -- 
    ra_14857_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => SHL_u32_u32_3776_inst_ack_0, ack => cp_elements(1106)); -- 
    -- CP-element group 1107 transition  input  bypass 
    -- predecessors 1104 
    -- successors 1112 
    -- members (7) 
      -- 	branch_block_stmt_2042/assign_stmt_3777_to_assign_stmt_3788/SHL_u32_u32_3776_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3777_to_assign_stmt_3788/SHL_u32_u32_3776_Update/$exit
      -- 	branch_block_stmt_2042/assign_stmt_3777_to_assign_stmt_3788/SHL_u32_u32_3776_Update/ca
      -- 	branch_block_stmt_2042/assign_stmt_3777_to_assign_stmt_3788/R_iNsTr_234_3785_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_3777_to_assign_stmt_3788/R_iNsTr_234_3785_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3777_to_assign_stmt_3788/R_iNsTr_234_3785_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_3777_to_assign_stmt_3788/R_iNsTr_234_3785_update_completed_
      -- 
    ca_14862_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => SHL_u32_u32_3776_inst_ack_1, ack => cp_elements(1107)); -- 
    -- CP-element group 1108 transition  output  bypass 
    -- predecessors 1103 
    -- successors 1111 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_3777_to_assign_stmt_3788/SHL_u32_u32_3782_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_3777_to_assign_stmt_3788/SHL_u32_u32_3782_Update/$entry
      -- 	branch_block_stmt_2042/assign_stmt_3777_to_assign_stmt_3788/SHL_u32_u32_3782_Update/cr
      -- 
    cp_elements(1108) <= cp_elements(1103);
    cr_14879_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1108), ack => SHL_u32_u32_3782_inst_req_1); -- 
    -- CP-element group 1109 transition  output  bypass 
    -- predecessors 1103 
    -- successors 1110 
    -- members (7) 
      -- 	branch_block_stmt_2042/assign_stmt_3777_to_assign_stmt_3788/SHL_u32_u32_3782_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_3777_to_assign_stmt_3788/R_curr_quotientx_x02x_xix_xi_3779_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_3777_to_assign_stmt_3788/R_curr_quotientx_x02x_xix_xi_3779_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3777_to_assign_stmt_3788/R_curr_quotientx_x02x_xix_xi_3779_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_3777_to_assign_stmt_3788/R_curr_quotientx_x02x_xix_xi_3779_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3777_to_assign_stmt_3788/SHL_u32_u32_3782_Sample/$entry
      -- 	branch_block_stmt_2042/assign_stmt_3777_to_assign_stmt_3788/SHL_u32_u32_3782_Sample/rr
      -- 
    cp_elements(1109) <= cp_elements(1103);
    rr_14874_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1109), ack => SHL_u32_u32_3782_inst_req_0); -- 
    -- CP-element group 1110 transition  input  bypass 
    -- predecessors 1109 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_3777_to_assign_stmt_3788/SHL_u32_u32_3782_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3777_to_assign_stmt_3788/SHL_u32_u32_3782_Sample/$exit
      -- 	branch_block_stmt_2042/assign_stmt_3777_to_assign_stmt_3788/SHL_u32_u32_3782_Sample/ra
      -- 
    ra_14875_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => SHL_u32_u32_3782_inst_ack_0, ack => cp_elements(1110)); -- 
    -- CP-element group 1111 transition  input  bypass 
    -- predecessors 1108 
    -- successors 1117 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_3777_to_assign_stmt_3788/SHL_u32_u32_3782_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3777_to_assign_stmt_3788/SHL_u32_u32_3782_Update/$exit
      -- 	branch_block_stmt_2042/assign_stmt_3777_to_assign_stmt_3788/SHL_u32_u32_3782_Update/ca
      -- 
    ca_14880_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => SHL_u32_u32_3782_inst_ack_1, ack => cp_elements(1111)); -- 
    -- CP-element group 1112 join  transition  output  bypass 
    -- predecessors 1107 1114 
    -- successors 1115 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_3777_to_assign_stmt_3788/ULT_u32_u1_3787_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_3777_to_assign_stmt_3788/ULT_u32_u1_3787_Sample/$entry
      -- 	branch_block_stmt_2042/assign_stmt_3777_to_assign_stmt_3788/ULT_u32_u1_3787_Sample/rr
      -- 
    cp_element_group_1112: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1112"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1107) & cp_elements(1114);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1112), clk => clk, reset => reset); --
    end block;
    rr_14896_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1112), ack => ULT_u32_u1_3787_inst_req_0); -- 
    -- CP-element group 1113 transition  output  bypass 
    -- predecessors 1103 
    -- successors 1116 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_3777_to_assign_stmt_3788/ULT_u32_u1_3787_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_3777_to_assign_stmt_3788/ULT_u32_u1_3787_Update/$entry
      -- 	branch_block_stmt_2042/assign_stmt_3777_to_assign_stmt_3788/ULT_u32_u1_3787_Update/cr
      -- 
    cp_elements(1113) <= cp_elements(1103);
    cr_14901_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1113), ack => ULT_u32_u1_3787_inst_req_1); -- 
    -- CP-element group 1114 transition  bypass 
    -- predecessors 1103 
    -- successors 1112 
    -- members (4) 
      -- 	branch_block_stmt_2042/assign_stmt_3777_to_assign_stmt_3788/R_iNsTr_183_3786_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_3777_to_assign_stmt_3788/R_iNsTr_183_3786_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3777_to_assign_stmt_3788/R_iNsTr_183_3786_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_3777_to_assign_stmt_3788/R_iNsTr_183_3786_update_completed_
      -- 
    cp_elements(1114) <= cp_elements(1103);
    -- CP-element group 1115 transition  input  bypass 
    -- predecessors 1112 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_3777_to_assign_stmt_3788/ULT_u32_u1_3787_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3777_to_assign_stmt_3788/ULT_u32_u1_3787_Sample/$exit
      -- 	branch_block_stmt_2042/assign_stmt_3777_to_assign_stmt_3788/ULT_u32_u1_3787_Sample/ra
      -- 
    ra_14897_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ULT_u32_u1_3787_inst_ack_0, ack => cp_elements(1115)); -- 
    -- CP-element group 1116 transition  input  bypass 
    -- predecessors 1113 
    -- successors 1117 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_3777_to_assign_stmt_3788/ULT_u32_u1_3787_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3777_to_assign_stmt_3788/ULT_u32_u1_3787_Update/$exit
      -- 	branch_block_stmt_2042/assign_stmt_3777_to_assign_stmt_3788/ULT_u32_u1_3787_Update/ca
      -- 
    ca_14902_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ULT_u32_u1_3787_inst_ack_1, ack => cp_elements(1116)); -- 
    -- CP-element group 1117 join  transition  bypass 
    -- predecessors 1111 1116 
    -- successors 68 
    -- members (1) 
      -- 	branch_block_stmt_2042/assign_stmt_3777_to_assign_stmt_3788/$exit
      -- 
    cp_element_group_1117: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1117"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1111) & cp_elements(1116);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1117), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1118 transition  place  dead  bypass 
    -- predecessors 68 
    -- successors 69 
    -- members (8) 
      -- 	branch_block_stmt_2042/if_stmt_3789__exit__
      -- 	branch_block_stmt_2042/merge_stmt_3795__entry__
      -- 	branch_block_stmt_2042/if_stmt_3789_dead_link/$entry
      -- 	branch_block_stmt_2042/if_stmt_3789_dead_link/$exit
      -- 	branch_block_stmt_2042/if_stmt_3789_dead_link/dead_transition
      -- 	branch_block_stmt_2042/merge_stmt_3795_dead_link/$entry
      -- 	branch_block_stmt_2042/merge_stmt_3795_dead_link/$exit
      -- 	branch_block_stmt_2042/merge_stmt_3795_dead_link/dead_transition
      -- 
    cp_elements(1118) <= false;
    -- CP-element group 1119 transition  output  bypass 
    -- predecessors 68 
    -- successors 1120 
    -- members (3) 
      -- 	branch_block_stmt_2042/if_stmt_3789_eval_test/$entry
      -- 	branch_block_stmt_2042/if_stmt_3789_eval_test/$exit
      -- 	branch_block_stmt_2042/if_stmt_3789_eval_test/branch_req
      -- 
    cp_elements(1119) <= cp_elements(68);
    branch_req_14910_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1119), ack => if_stmt_3789_branch_req_0); -- 
    -- CP-element group 1120 branch  place  bypass 
    -- predecessors 1119 
    -- successors 1121 1123 
    -- members (1) 
      -- 	branch_block_stmt_2042/R_iNsTr_236_3790_place
      -- 
    cp_elements(1120) <= cp_elements(1119);
    -- CP-element group 1121 transition  bypass 
    -- predecessors 1120 
    -- successors 1122 
    -- members (1) 
      -- 	branch_block_stmt_2042/if_stmt_3789_if_link/$entry
      -- 
    cp_elements(1121) <= cp_elements(1120);
    -- CP-element group 1122 transition  place  input  bypass 
    -- predecessors 1121 
    -- successors 2373 
    -- members (3) 
      -- 	branch_block_stmt_2042/if_stmt_3789_if_link/$exit
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xi_bbx_xnphx_xix_xi
      -- 	branch_block_stmt_2042/if_stmt_3789_if_link/if_choice_transition
      -- 
    if_choice_transition_14915_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_3789_branch_ack_1, ack => cp_elements(1122)); -- 
    -- CP-element group 1123 transition  bypass 
    -- predecessors 1120 
    -- successors 1124 
    -- members (1) 
      -- 	branch_block_stmt_2042/if_stmt_3789_else_link/$entry
      -- 
    cp_elements(1123) <= cp_elements(1120);
    -- CP-element group 1124 transition  place  input  bypass 
    -- predecessors 1123 
    -- successors 2402 
    -- members (3) 
      -- 	branch_block_stmt_2042/if_stmt_3789_else_link/$exit
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xi_xx_x_crit_edgex_xix_xix_xloopexit
      -- 	branch_block_stmt_2042/if_stmt_3789_else_link/else_choice_transition
      -- 
    else_choice_transition_14919_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_3789_branch_ack_0, ack => cp_elements(1124)); -- 
    -- CP-element group 1125 fork  transition  bypass 
    -- predecessors 70 
    -- successors 1127 1128 1129 1133 1134 1135 1138 
    -- members (1) 
      -- 	branch_block_stmt_2042/assign_stmt_3826_to_assign_stmt_3837/$entry
      -- 
    cp_elements(1125) <= cp_elements(70);
    -- CP-element group 1126 join  transition  output  bypass 
    -- predecessors 1128 1129 
    -- successors 1130 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_3826_to_assign_stmt_3837/ADD_u32_u32_3825_Sample/$entry
      -- 	branch_block_stmt_2042/assign_stmt_3826_to_assign_stmt_3837/ADD_u32_u32_3825_Sample/rr
      -- 	branch_block_stmt_2042/assign_stmt_3826_to_assign_stmt_3837/ADD_u32_u32_3825_sample_start_
      -- 
    cp_element_group_1126: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1126"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1128) & cp_elements(1129);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1126), clk => clk, reset => reset); --
    end block;
    rr_14940_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1126), ack => ADD_u32_u32_3825_inst_req_0); -- 
    -- CP-element group 1127 transition  output  bypass 
    -- predecessors 1125 
    -- successors 1131 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_3826_to_assign_stmt_3837/ADD_u32_u32_3825_Update/$entry
      -- 	branch_block_stmt_2042/assign_stmt_3826_to_assign_stmt_3837/ADD_u32_u32_3825_Update/cr
      -- 	branch_block_stmt_2042/assign_stmt_3826_to_assign_stmt_3837/ADD_u32_u32_3825_update_start_
      -- 
    cp_elements(1127) <= cp_elements(1125);
    cr_14945_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1127), ack => ADD_u32_u32_3825_inst_req_1); -- 
    -- CP-element group 1128 transition  bypass 
    -- predecessors 1125 
    -- successors 1126 
    -- members (4) 
      -- 	branch_block_stmt_2042/assign_stmt_3826_to_assign_stmt_3837/R_curr_quotientx_x0x_xlcssax_xix_xi_3823_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3826_to_assign_stmt_3837/R_curr_quotientx_x0x_xlcssax_xix_xi_3823_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_3826_to_assign_stmt_3837/R_curr_quotientx_x0x_xlcssax_xix_xi_3823_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3826_to_assign_stmt_3837/R_curr_quotientx_x0x_xlcssax_xix_xi_3823_sample_start_
      -- 
    cp_elements(1128) <= cp_elements(1125);
    -- CP-element group 1129 transition  bypass 
    -- predecessors 1125 
    -- successors 1126 
    -- members (4) 
      -- 	branch_block_stmt_2042/assign_stmt_3826_to_assign_stmt_3837/R_quotientx_x05x_xix_xi_3824_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_3826_to_assign_stmt_3837/R_quotientx_x05x_xix_xi_3824_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3826_to_assign_stmt_3837/R_quotientx_x05x_xix_xi_3824_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_3826_to_assign_stmt_3837/R_quotientx_x05x_xix_xi_3824_sample_completed_
      -- 
    cp_elements(1129) <= cp_elements(1125);
    -- CP-element group 1130 transition  input  bypass 
    -- predecessors 1126 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_3826_to_assign_stmt_3837/ADD_u32_u32_3825_Sample/$exit
      -- 	branch_block_stmt_2042/assign_stmt_3826_to_assign_stmt_3837/ADD_u32_u32_3825_Sample/ra
      -- 	branch_block_stmt_2042/assign_stmt_3826_to_assign_stmt_3837/ADD_u32_u32_3825_sample_completed_
      -- 
    ra_14941_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u32_u32_3825_inst_ack_0, ack => cp_elements(1130)); -- 
    -- CP-element group 1131 transition  input  bypass 
    -- predecessors 1127 
    -- successors 1141 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_3826_to_assign_stmt_3837/ADD_u32_u32_3825_Update/$exit
      -- 	branch_block_stmt_2042/assign_stmt_3826_to_assign_stmt_3837/ADD_u32_u32_3825_Update/ca
      -- 	branch_block_stmt_2042/assign_stmt_3826_to_assign_stmt_3837/ADD_u32_u32_3825_update_completed_
      -- 
    ca_14946_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u32_u32_3825_inst_ack_1, ack => cp_elements(1131)); -- 
    -- CP-element group 1132 join  transition  output  bypass 
    -- predecessors 1134 1135 
    -- successors 1136 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_3826_to_assign_stmt_3837/SUB_u32_u32_3830_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_3826_to_assign_stmt_3837/SUB_u32_u32_3830_Sample/rr
      -- 	branch_block_stmt_2042/assign_stmt_3826_to_assign_stmt_3837/SUB_u32_u32_3830_Sample/$entry
      -- 
    cp_element_group_1132: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1132"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1134) & cp_elements(1135);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1132), clk => clk, reset => reset); --
    end block;
    rr_14962_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1132), ack => SUB_u32_u32_3830_inst_req_0); -- 
    -- CP-element group 1133 transition  output  bypass 
    -- predecessors 1125 
    -- successors 1137 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_3826_to_assign_stmt_3837/SUB_u32_u32_3830_Update/cr
      -- 	branch_block_stmt_2042/assign_stmt_3826_to_assign_stmt_3837/SUB_u32_u32_3830_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_3826_to_assign_stmt_3837/SUB_u32_u32_3830_Update/$entry
      -- 
    cp_elements(1133) <= cp_elements(1125);
    cr_14967_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1133), ack => SUB_u32_u32_3830_inst_req_1); -- 
    -- CP-element group 1134 transition  bypass 
    -- predecessors 1125 
    -- successors 1132 
    -- members (4) 
      -- 	branch_block_stmt_2042/assign_stmt_3826_to_assign_stmt_3837/R_xx_x016x_xix_xi_3828_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_3826_to_assign_stmt_3837/R_xx_x016x_xix_xi_3828_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3826_to_assign_stmt_3837/R_xx_x016x_xix_xi_3828_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_3826_to_assign_stmt_3837/R_xx_x016x_xix_xi_3828_update_completed_
      -- 
    cp_elements(1134) <= cp_elements(1125);
    -- CP-element group 1135 transition  bypass 
    -- predecessors 1125 
    -- successors 1132 
    -- members (4) 
      -- 	branch_block_stmt_2042/assign_stmt_3826_to_assign_stmt_3837/R_shifted_divisorx_x0x_xlcssax_xix_xi_3829_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_3826_to_assign_stmt_3837/R_shifted_divisorx_x0x_xlcssax_xix_xi_3829_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3826_to_assign_stmt_3837/R_shifted_divisorx_x0x_xlcssax_xix_xi_3829_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_3826_to_assign_stmt_3837/R_shifted_divisorx_x0x_xlcssax_xix_xi_3829_update_completed_
      -- 
    cp_elements(1135) <= cp_elements(1125);
    -- CP-element group 1136 transition  input  bypass 
    -- predecessors 1132 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_3826_to_assign_stmt_3837/SUB_u32_u32_3830_Sample/$exit
      -- 	branch_block_stmt_2042/assign_stmt_3826_to_assign_stmt_3837/SUB_u32_u32_3830_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3826_to_assign_stmt_3837/SUB_u32_u32_3830_Sample/ra
      -- 
    ra_14963_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => SUB_u32_u32_3830_inst_ack_0, ack => cp_elements(1136)); -- 
    -- CP-element group 1137 transition  input  output  bypass 
    -- predecessors 1133 
    -- successors 1139 
    -- members (10) 
      -- 	branch_block_stmt_2042/assign_stmt_3826_to_assign_stmt_3837/SUB_u32_u32_3830_Update/$exit
      -- 	branch_block_stmt_2042/assign_stmt_3826_to_assign_stmt_3837/R_iNsTr_213_3833_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_3826_to_assign_stmt_3837/R_iNsTr_213_3833_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3826_to_assign_stmt_3837/R_iNsTr_213_3833_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_3826_to_assign_stmt_3837/R_iNsTr_213_3833_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3826_to_assign_stmt_3837/ULT_u32_u1_3836_Sample/$entry
      -- 	branch_block_stmt_2042/assign_stmt_3826_to_assign_stmt_3837/SUB_u32_u32_3830_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3826_to_assign_stmt_3837/ULT_u32_u1_3836_Sample/rr
      -- 	branch_block_stmt_2042/assign_stmt_3826_to_assign_stmt_3837/ULT_u32_u1_3836_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_3826_to_assign_stmt_3837/SUB_u32_u32_3830_Update/ca
      -- 
    ca_14968_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => SUB_u32_u32_3830_inst_ack_1, ack => cp_elements(1137)); -- 
    rr_14980_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1137), ack => ULT_u32_u1_3836_inst_req_0); -- 
    -- CP-element group 1138 transition  output  bypass 
    -- predecessors 1125 
    -- successors 1140 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_3826_to_assign_stmt_3837/ULT_u32_u1_3836_Update/$entry
      -- 	branch_block_stmt_2042/assign_stmt_3826_to_assign_stmt_3837/ULT_u32_u1_3836_Update/cr
      -- 	branch_block_stmt_2042/assign_stmt_3826_to_assign_stmt_3837/ULT_u32_u1_3836_update_start_
      -- 
    cp_elements(1138) <= cp_elements(1125);
    cr_14985_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1138), ack => ULT_u32_u1_3836_inst_req_1); -- 
    -- CP-element group 1139 transition  input  bypass 
    -- predecessors 1137 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_3826_to_assign_stmt_3837/ULT_u32_u1_3836_Sample/$exit
      -- 	branch_block_stmt_2042/assign_stmt_3826_to_assign_stmt_3837/ULT_u32_u1_3836_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3826_to_assign_stmt_3837/ULT_u32_u1_3836_Sample/ra
      -- 
    ra_14981_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ULT_u32_u1_3836_inst_ack_0, ack => cp_elements(1139)); -- 
    -- CP-element group 1140 transition  input  bypass 
    -- predecessors 1138 
    -- successors 1141 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_3826_to_assign_stmt_3837/ULT_u32_u1_3836_Update/$exit
      -- 	branch_block_stmt_2042/assign_stmt_3826_to_assign_stmt_3837/ULT_u32_u1_3836_Update/ca
      -- 	branch_block_stmt_2042/assign_stmt_3826_to_assign_stmt_3837/ULT_u32_u1_3836_update_completed_
      -- 
    ca_14986_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ULT_u32_u1_3836_inst_ack_1, ack => cp_elements(1140)); -- 
    -- CP-element group 1141 join  transition  bypass 
    -- predecessors 1131 1140 
    -- successors 71 
    -- members (1) 
      -- 	branch_block_stmt_2042/assign_stmt_3826_to_assign_stmt_3837/$exit
      -- 
    cp_element_group_1141: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1141"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1131) & cp_elements(1140);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1141), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1142 transition  place  dead  bypass 
    -- predecessors 71 
    -- successors 72 
    -- members (8) 
      -- 	branch_block_stmt_2042/if_stmt_3838__exit__
      -- 	branch_block_stmt_2042/merge_stmt_3844__entry__
      -- 	branch_block_stmt_2042/if_stmt_3838_dead_link/dead_transition
      -- 	branch_block_stmt_2042/if_stmt_3838_dead_link/$entry
      -- 	branch_block_stmt_2042/if_stmt_3838_dead_link/$exit
      -- 	branch_block_stmt_2042/merge_stmt_3844_dead_link/$entry
      -- 	branch_block_stmt_2042/merge_stmt_3844_dead_link/$exit
      -- 	branch_block_stmt_2042/merge_stmt_3844_dead_link/dead_transition
      -- 
    cp_elements(1142) <= false;
    -- CP-element group 1143 transition  output  bypass 
    -- predecessors 71 
    -- successors 1144 
    -- members (3) 
      -- 	branch_block_stmt_2042/if_stmt_3838_eval_test/$entry
      -- 	branch_block_stmt_2042/if_stmt_3838_eval_test/$exit
      -- 	branch_block_stmt_2042/if_stmt_3838_eval_test/branch_req
      -- 
    cp_elements(1143) <= cp_elements(71);
    branch_req_14994_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1143), ack => if_stmt_3838_branch_req_0); -- 
    -- CP-element group 1144 branch  place  bypass 
    -- predecessors 1143 
    -- successors 1145 1147 
    -- members (1) 
      -- 	branch_block_stmt_2042/R_iNsTr_214_3839_place
      -- 
    cp_elements(1144) <= cp_elements(1143);
    -- CP-element group 1145 transition  bypass 
    -- predecessors 1144 
    -- successors 1146 
    -- members (1) 
      -- 	branch_block_stmt_2042/if_stmt_3838_if_link/$entry
      -- 
    cp_elements(1145) <= cp_elements(1144);
    -- CP-element group 1146 fork  transition  place  input  bypass 
    -- predecessors 1145 
    -- successors 2450 2452 
    -- members (8) 
      -- 	branch_block_stmt_2042/if_stmt_3838_if_link/if_choice_transition
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xi_udiv32x_xexitx_xpreheaderx_xi
      -- 	branch_block_stmt_2042/if_stmt_3838_if_link/$exit
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xi_udiv32x_xexitx_xpreheaderx_xi_PhiReq/$entry
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xi_udiv32x_xexitx_xpreheaderx_xi_PhiReq/phi_stmt_3845/$entry
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xi_udiv32x_xexitx_xpreheaderx_xi_PhiReq/phi_stmt_3845/phi_stmt_3845_sources/$entry
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xi_udiv32x_xexitx_xpreheaderx_xi_PhiReq/phi_stmt_3845/phi_stmt_3845_sources/type_cast_3848/$entry
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xi_udiv32x_xexitx_xpreheaderx_xi_PhiReq/phi_stmt_3845/phi_stmt_3845_sources/type_cast_3848/SplitProtocol/$entry
      -- 
    if_choice_transition_14999_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_3838_branch_ack_1, ack => cp_elements(1146)); -- 
    -- CP-element group 1147 transition  bypass 
    -- predecessors 1144 
    -- successors 1148 
    -- members (1) 
      -- 	branch_block_stmt_2042/if_stmt_3838_else_link/$entry
      -- 
    cp_elements(1147) <= cp_elements(1144);
    -- CP-element group 1148 transition  place  input  bypass 
    -- predecessors 1147 
    -- successors 2330 
    -- members (3) 
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xi_bbx_xnph7x_xix_xi
      -- 	branch_block_stmt_2042/if_stmt_3838_else_link/$exit
      -- 	branch_block_stmt_2042/if_stmt_3838_else_link/else_choice_transition
      -- 
    else_choice_transition_15003_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_3838_branch_ack_0, ack => cp_elements(1148)); -- 
    -- CP-element group 1149 fork  transition  bypass 
    -- predecessors 72 
    -- successors 1150 1151 1154 1155 1158 1161 1164 1165 1168 1171 1172 1178 
    -- members (1) 
      -- 	branch_block_stmt_2042/assign_stmt_3855_to_assign_stmt_3898/$entry
      -- 
    cp_elements(1149) <= cp_elements(72);
    -- CP-element group 1150 transition  output  bypass 
    -- predecessors 1149 
    -- successors 1153 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_3855_to_assign_stmt_3898/LSHR_u32_u32_3854_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_3855_to_assign_stmt_3898/LSHR_u32_u32_3854_Update/$entry
      -- 	branch_block_stmt_2042/assign_stmt_3855_to_assign_stmt_3898/LSHR_u32_u32_3854_Update/cr
      -- 
    cp_elements(1150) <= cp_elements(1149);
    cr_15025_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1150), ack => LSHR_u32_u32_3854_inst_req_1); -- 
    -- CP-element group 1151 transition  output  bypass 
    -- predecessors 1149 
    -- successors 1152 
    -- members (7) 
      -- 	branch_block_stmt_2042/assign_stmt_3855_to_assign_stmt_3898/LSHR_u32_u32_3854_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_3855_to_assign_stmt_3898/R_tmp10x_xi55_3851_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_3855_to_assign_stmt_3898/R_tmp10x_xi55_3851_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3855_to_assign_stmt_3898/R_tmp10x_xi55_3851_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_3855_to_assign_stmt_3898/R_tmp10x_xi55_3851_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3855_to_assign_stmt_3898/LSHR_u32_u32_3854_Sample/$entry
      -- 	branch_block_stmt_2042/assign_stmt_3855_to_assign_stmt_3898/LSHR_u32_u32_3854_Sample/rr
      -- 
    cp_elements(1151) <= cp_elements(1149);
    rr_15020_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1151), ack => LSHR_u32_u32_3854_inst_req_0); -- 
    -- CP-element group 1152 transition  input  bypass 
    -- predecessors 1151 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_3855_to_assign_stmt_3898/LSHR_u32_u32_3854_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3855_to_assign_stmt_3898/LSHR_u32_u32_3854_Sample/$exit
      -- 	branch_block_stmt_2042/assign_stmt_3855_to_assign_stmt_3898/LSHR_u32_u32_3854_Sample/ra
      -- 
    ra_15021_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => LSHR_u32_u32_3854_inst_ack_0, ack => cp_elements(1152)); -- 
    -- CP-element group 1153 transition  input  output  bypass 
    -- predecessors 1150 
    -- successors 1159 
    -- members (10) 
      -- 	branch_block_stmt_2042/assign_stmt_3855_to_assign_stmt_3898/LSHR_u32_u32_3854_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3855_to_assign_stmt_3898/LSHR_u32_u32_3854_Update/$exit
      -- 	branch_block_stmt_2042/assign_stmt_3855_to_assign_stmt_3898/LSHR_u32_u32_3854_Update/ca
      -- 	branch_block_stmt_2042/assign_stmt_3855_to_assign_stmt_3898/AND_u32_u32_3866_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_3855_to_assign_stmt_3898/R_iNsTr_238_3863_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_3855_to_assign_stmt_3898/R_iNsTr_238_3863_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3855_to_assign_stmt_3898/R_iNsTr_238_3863_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_3855_to_assign_stmt_3898/R_iNsTr_238_3863_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3855_to_assign_stmt_3898/AND_u32_u32_3866_Sample/$entry
      -- 	branch_block_stmt_2042/assign_stmt_3855_to_assign_stmt_3898/AND_u32_u32_3866_Sample/rr
      -- 
    ca_15026_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => LSHR_u32_u32_3854_inst_ack_1, ack => cp_elements(1153)); -- 
    rr_15056_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1153), ack => AND_u32_u32_3866_inst_req_0); -- 
    -- CP-element group 1154 transition  output  bypass 
    -- predecessors 1149 
    -- successors 1157 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_3855_to_assign_stmt_3898/AND_u32_u32_3860_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_3855_to_assign_stmt_3898/AND_u32_u32_3860_Update/$entry
      -- 	branch_block_stmt_2042/assign_stmt_3855_to_assign_stmt_3898/AND_u32_u32_3860_Update/cr
      -- 
    cp_elements(1154) <= cp_elements(1149);
    cr_15043_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1154), ack => AND_u32_u32_3860_inst_req_1); -- 
    -- CP-element group 1155 transition  output  bypass 
    -- predecessors 1149 
    -- successors 1156 
    -- members (7) 
      -- 	branch_block_stmt_2042/assign_stmt_3855_to_assign_stmt_3898/AND_u32_u32_3860_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_3855_to_assign_stmt_3898/R_tmp10x_xi55_3857_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_3855_to_assign_stmt_3898/R_tmp10x_xi55_3857_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3855_to_assign_stmt_3898/R_tmp10x_xi55_3857_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_3855_to_assign_stmt_3898/R_tmp10x_xi55_3857_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3855_to_assign_stmt_3898/AND_u32_u32_3860_Sample/$entry
      -- 	branch_block_stmt_2042/assign_stmt_3855_to_assign_stmt_3898/AND_u32_u32_3860_Sample/rr
      -- 
    cp_elements(1155) <= cp_elements(1149);
    rr_15038_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1155), ack => AND_u32_u32_3860_inst_req_0); -- 
    -- CP-element group 1156 transition  input  bypass 
    -- predecessors 1155 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_3855_to_assign_stmt_3898/AND_u32_u32_3860_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3855_to_assign_stmt_3898/AND_u32_u32_3860_Sample/$exit
      -- 	branch_block_stmt_2042/assign_stmt_3855_to_assign_stmt_3898/AND_u32_u32_3860_Sample/ra
      -- 
    ra_15039_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => AND_u32_u32_3860_inst_ack_0, ack => cp_elements(1156)); -- 
    -- CP-element group 1157 transition  input  bypass 
    -- predecessors 1154 
    -- successors 1181 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_3855_to_assign_stmt_3898/AND_u32_u32_3860_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3855_to_assign_stmt_3898/AND_u32_u32_3860_Update/$exit
      -- 	branch_block_stmt_2042/assign_stmt_3855_to_assign_stmt_3898/AND_u32_u32_3860_Update/ca
      -- 
    ca_15044_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => AND_u32_u32_3860_inst_ack_1, ack => cp_elements(1157)); -- 
    -- CP-element group 1158 transition  output  bypass 
    -- predecessors 1149 
    -- successors 1160 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_3855_to_assign_stmt_3898/AND_u32_u32_3866_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_3855_to_assign_stmt_3898/AND_u32_u32_3866_Update/$entry
      -- 	branch_block_stmt_2042/assign_stmt_3855_to_assign_stmt_3898/AND_u32_u32_3866_Update/cr
      -- 
    cp_elements(1158) <= cp_elements(1149);
    cr_15061_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1158), ack => AND_u32_u32_3866_inst_req_1); -- 
    -- CP-element group 1159 transition  input  bypass 
    -- predecessors 1153 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_3855_to_assign_stmt_3898/AND_u32_u32_3866_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3855_to_assign_stmt_3898/AND_u32_u32_3866_Sample/$exit
      -- 	branch_block_stmt_2042/assign_stmt_3855_to_assign_stmt_3898/AND_u32_u32_3866_Sample/ra
      -- 
    ra_15057_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => AND_u32_u32_3866_inst_ack_0, ack => cp_elements(1159)); -- 
    -- CP-element group 1160 transition  input  output  bypass 
    -- predecessors 1158 
    -- successors 1162 
    -- members (10) 
      -- 	branch_block_stmt_2042/assign_stmt_3855_to_assign_stmt_3898/AND_u32_u32_3866_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3855_to_assign_stmt_3898/AND_u32_u32_3866_Update/$exit
      -- 	branch_block_stmt_2042/assign_stmt_3855_to_assign_stmt_3898/AND_u32_u32_3866_Update/ca
      -- 	branch_block_stmt_2042/assign_stmt_3855_to_assign_stmt_3898/ADD_u32_u32_3872_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_3855_to_assign_stmt_3898/R_iNsTr_240_3869_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_3855_to_assign_stmt_3898/R_iNsTr_240_3869_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3855_to_assign_stmt_3898/R_iNsTr_240_3869_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_3855_to_assign_stmt_3898/R_iNsTr_240_3869_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3855_to_assign_stmt_3898/ADD_u32_u32_3872_Sample/$entry
      -- 	branch_block_stmt_2042/assign_stmt_3855_to_assign_stmt_3898/ADD_u32_u32_3872_Sample/rr
      -- 
    ca_15062_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => AND_u32_u32_3866_inst_ack_1, ack => cp_elements(1160)); -- 
    rr_15074_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1160), ack => ADD_u32_u32_3872_inst_req_0); -- 
    -- CP-element group 1161 transition  output  bypass 
    -- predecessors 1149 
    -- successors 1163 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_3855_to_assign_stmt_3898/ADD_u32_u32_3872_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_3855_to_assign_stmt_3898/ADD_u32_u32_3872_Update/$entry
      -- 	branch_block_stmt_2042/assign_stmt_3855_to_assign_stmt_3898/ADD_u32_u32_3872_Update/cr
      -- 
    cp_elements(1161) <= cp_elements(1149);
    cr_15079_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1161), ack => ADD_u32_u32_3872_inst_req_1); -- 
    -- CP-element group 1162 transition  input  bypass 
    -- predecessors 1160 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_3855_to_assign_stmt_3898/ADD_u32_u32_3872_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3855_to_assign_stmt_3898/ADD_u32_u32_3872_Sample/$exit
      -- 	branch_block_stmt_2042/assign_stmt_3855_to_assign_stmt_3898/ADD_u32_u32_3872_Sample/ra
      -- 
    ra_15075_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u32_u32_3872_inst_ack_0, ack => cp_elements(1162)); -- 
    -- CP-element group 1163 transition  input  bypass 
    -- predecessors 1161 
    -- successors 1181 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_3855_to_assign_stmt_3898/ADD_u32_u32_3872_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3855_to_assign_stmt_3898/ADD_u32_u32_3872_Update/$exit
      -- 	branch_block_stmt_2042/assign_stmt_3855_to_assign_stmt_3898/ADD_u32_u32_3872_Update/ca
      -- 
    ca_15080_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u32_u32_3872_inst_ack_1, ack => cp_elements(1163)); -- 
    -- CP-element group 1164 transition  output  bypass 
    -- predecessors 1149 
    -- successors 1167 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_3855_to_assign_stmt_3898/AND_u32_u32_3878_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_3855_to_assign_stmt_3898/AND_u32_u32_3878_Update/$entry
      -- 	branch_block_stmt_2042/assign_stmt_3855_to_assign_stmt_3898/AND_u32_u32_3878_Update/cr
      -- 
    cp_elements(1164) <= cp_elements(1149);
    cr_15097_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1164), ack => AND_u32_u32_3878_inst_req_1); -- 
    -- CP-element group 1165 transition  output  bypass 
    -- predecessors 1149 
    -- successors 1166 
    -- members (7) 
      -- 	branch_block_stmt_2042/assign_stmt_3855_to_assign_stmt_3898/AND_u32_u32_3878_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_3855_to_assign_stmt_3898/R_xx_xlcssa4_3875_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_3855_to_assign_stmt_3898/R_xx_xlcssa4_3875_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3855_to_assign_stmt_3898/R_xx_xlcssa4_3875_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_3855_to_assign_stmt_3898/R_xx_xlcssa4_3875_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3855_to_assign_stmt_3898/AND_u32_u32_3878_Sample/$entry
      -- 	branch_block_stmt_2042/assign_stmt_3855_to_assign_stmt_3898/AND_u32_u32_3878_Sample/rr
      -- 
    cp_elements(1165) <= cp_elements(1149);
    rr_15092_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1165), ack => AND_u32_u32_3878_inst_req_0); -- 
    -- CP-element group 1166 transition  input  bypass 
    -- predecessors 1165 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_3855_to_assign_stmt_3898/AND_u32_u32_3878_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3855_to_assign_stmt_3898/AND_u32_u32_3878_Sample/$exit
      -- 	branch_block_stmt_2042/assign_stmt_3855_to_assign_stmt_3898/AND_u32_u32_3878_Sample/ra
      -- 
    ra_15093_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => AND_u32_u32_3878_inst_ack_0, ack => cp_elements(1166)); -- 
    -- CP-element group 1167 transition  input  output  bypass 
    -- predecessors 1164 
    -- successors 1169 
    -- members (10) 
      -- 	branch_block_stmt_2042/assign_stmt_3855_to_assign_stmt_3898/AND_u32_u32_3878_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3855_to_assign_stmt_3898/AND_u32_u32_3878_Update/$exit
      -- 	branch_block_stmt_2042/assign_stmt_3855_to_assign_stmt_3898/AND_u32_u32_3878_Update/ca
      -- 	branch_block_stmt_2042/assign_stmt_3855_to_assign_stmt_3898/EQ_u32_u1_3884_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_3855_to_assign_stmt_3898/R_iNsTr_242_3881_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_3855_to_assign_stmt_3898/R_iNsTr_242_3881_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3855_to_assign_stmt_3898/R_iNsTr_242_3881_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_3855_to_assign_stmt_3898/R_iNsTr_242_3881_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3855_to_assign_stmt_3898/EQ_u32_u1_3884_Sample/$entry
      -- 	branch_block_stmt_2042/assign_stmt_3855_to_assign_stmt_3898/EQ_u32_u1_3884_Sample/rr
      -- 
    ca_15098_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => AND_u32_u32_3878_inst_ack_1, ack => cp_elements(1167)); -- 
    rr_15110_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1167), ack => EQ_u32_u1_3884_inst_req_0); -- 
    -- CP-element group 1168 transition  output  bypass 
    -- predecessors 1149 
    -- successors 1170 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_3855_to_assign_stmt_3898/EQ_u32_u1_3884_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_3855_to_assign_stmt_3898/EQ_u32_u1_3884_Update/$entry
      -- 	branch_block_stmt_2042/assign_stmt_3855_to_assign_stmt_3898/EQ_u32_u1_3884_Update/cr
      -- 
    cp_elements(1168) <= cp_elements(1149);
    cr_15115_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1168), ack => EQ_u32_u1_3884_inst_req_1); -- 
    -- CP-element group 1169 transition  input  bypass 
    -- predecessors 1167 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_3855_to_assign_stmt_3898/EQ_u32_u1_3884_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3855_to_assign_stmt_3898/EQ_u32_u1_3884_Sample/$exit
      -- 	branch_block_stmt_2042/assign_stmt_3855_to_assign_stmt_3898/EQ_u32_u1_3884_Sample/ra
      -- 
    ra_15111_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u32_u1_3884_inst_ack_0, ack => cp_elements(1169)); -- 
    -- CP-element group 1170 transition  input  bypass 
    -- predecessors 1168 
    -- successors 1177 
    -- members (7) 
      -- 	branch_block_stmt_2042/assign_stmt_3855_to_assign_stmt_3898/EQ_u32_u1_3884_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3855_to_assign_stmt_3898/EQ_u32_u1_3884_Update/$exit
      -- 	branch_block_stmt_2042/assign_stmt_3855_to_assign_stmt_3898/EQ_u32_u1_3884_Update/ca
      -- 	branch_block_stmt_2042/assign_stmt_3855_to_assign_stmt_3898/R_iNsTr_243_3895_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_3855_to_assign_stmt_3898/R_iNsTr_243_3895_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3855_to_assign_stmt_3898/R_iNsTr_243_3895_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_3855_to_assign_stmt_3898/R_iNsTr_243_3895_update_completed_
      -- 
    ca_15116_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u32_u1_3884_inst_ack_1, ack => cp_elements(1170)); -- 
    -- CP-element group 1171 transition  output  bypass 
    -- predecessors 1149 
    -- successors 1176 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_3855_to_assign_stmt_3898/NEQ_i32_u1_3892_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_3855_to_assign_stmt_3898/NEQ_i32_u1_3892_Update/$entry
      -- 	branch_block_stmt_2042/assign_stmt_3855_to_assign_stmt_3898/NEQ_i32_u1_3892_Update/cr
      -- 
    cp_elements(1171) <= cp_elements(1149);
    cr_15147_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1171), ack => NEQ_i32_u1_3892_inst_req_1); -- 
    -- CP-element group 1172 transition  output  bypass 
    -- predecessors 1149 
    -- successors 1173 
    -- members (7) 
      -- 	branch_block_stmt_2042/assign_stmt_3855_to_assign_stmt_3898/type_cast_3888_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_3855_to_assign_stmt_3898/R_xx_xlcssa4_3887_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_3855_to_assign_stmt_3898/R_xx_xlcssa4_3887_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3855_to_assign_stmt_3898/R_xx_xlcssa4_3887_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_3855_to_assign_stmt_3898/R_xx_xlcssa4_3887_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3855_to_assign_stmt_3898/type_cast_3888_Sample/$entry
      -- 	branch_block_stmt_2042/assign_stmt_3855_to_assign_stmt_3898/type_cast_3888_Sample/rr
      -- 
    cp_elements(1172) <= cp_elements(1149);
    rr_15132_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1172), ack => type_cast_3888_inst_req_0); -- 
    -- CP-element group 1173 transition  input  output  bypass 
    -- predecessors 1172 
    -- successors 1174 
    -- members (6) 
      -- 	branch_block_stmt_2042/assign_stmt_3855_to_assign_stmt_3898/type_cast_3888_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3855_to_assign_stmt_3898/type_cast_3888_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_3855_to_assign_stmt_3898/type_cast_3888_Sample/$exit
      -- 	branch_block_stmt_2042/assign_stmt_3855_to_assign_stmt_3898/type_cast_3888_Sample/ra
      -- 	branch_block_stmt_2042/assign_stmt_3855_to_assign_stmt_3898/type_cast_3888_Update/$entry
      -- 	branch_block_stmt_2042/assign_stmt_3855_to_assign_stmt_3898/type_cast_3888_Update/cr
      -- 
    ra_15133_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3888_inst_ack_0, ack => cp_elements(1173)); -- 
    cr_15137_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1173), ack => type_cast_3888_inst_req_1); -- 
    -- CP-element group 1174 transition  input  output  bypass 
    -- predecessors 1173 
    -- successors 1175 
    -- members (6) 
      -- 	branch_block_stmt_2042/assign_stmt_3855_to_assign_stmt_3898/NEQ_i32_u1_3892_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_3855_to_assign_stmt_3898/type_cast_3888_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3855_to_assign_stmt_3898/type_cast_3888_Update/$exit
      -- 	branch_block_stmt_2042/assign_stmt_3855_to_assign_stmt_3898/type_cast_3888_Update/ca
      -- 	branch_block_stmt_2042/assign_stmt_3855_to_assign_stmt_3898/NEQ_i32_u1_3892_Sample/$entry
      -- 	branch_block_stmt_2042/assign_stmt_3855_to_assign_stmt_3898/NEQ_i32_u1_3892_Sample/rr
      -- 
    ca_15138_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3888_inst_ack_1, ack => cp_elements(1174)); -- 
    rr_15142_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1174), ack => NEQ_i32_u1_3892_inst_req_0); -- 
    -- CP-element group 1175 transition  input  bypass 
    -- predecessors 1174 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_3855_to_assign_stmt_3898/NEQ_i32_u1_3892_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3855_to_assign_stmt_3898/NEQ_i32_u1_3892_Sample/$exit
      -- 	branch_block_stmt_2042/assign_stmt_3855_to_assign_stmt_3898/NEQ_i32_u1_3892_Sample/ra
      -- 
    ra_15143_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => NEQ_i32_u1_3892_inst_ack_0, ack => cp_elements(1175)); -- 
    -- CP-element group 1176 transition  input  bypass 
    -- predecessors 1171 
    -- successors 1177 
    -- members (7) 
      -- 	branch_block_stmt_2042/assign_stmt_3855_to_assign_stmt_3898/NEQ_i32_u1_3892_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3855_to_assign_stmt_3898/NEQ_i32_u1_3892_Update/$exit
      -- 	branch_block_stmt_2042/assign_stmt_3855_to_assign_stmt_3898/NEQ_i32_u1_3892_Update/ca
      -- 	branch_block_stmt_2042/assign_stmt_3855_to_assign_stmt_3898/R_iNsTr_244_3896_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_3855_to_assign_stmt_3898/R_iNsTr_244_3896_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3855_to_assign_stmt_3898/R_iNsTr_244_3896_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_3855_to_assign_stmt_3898/R_iNsTr_244_3896_update_completed_
      -- 
    ca_15148_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => NEQ_i32_u1_3892_inst_ack_1, ack => cp_elements(1176)); -- 
    -- CP-element group 1177 join  transition  output  bypass 
    -- predecessors 1170 1176 
    -- successors 1179 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_3855_to_assign_stmt_3898/AND_u1_u1_3897_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_3855_to_assign_stmt_3898/AND_u1_u1_3897_Sample/$entry
      -- 	branch_block_stmt_2042/assign_stmt_3855_to_assign_stmt_3898/AND_u1_u1_3897_Sample/rr
      -- 
    cp_element_group_1177: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1177"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1170) & cp_elements(1176);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1177), clk => clk, reset => reset); --
    end block;
    rr_15164_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1177), ack => AND_u1_u1_3897_inst_req_0); -- 
    -- CP-element group 1178 transition  output  bypass 
    -- predecessors 1149 
    -- successors 1180 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_3855_to_assign_stmt_3898/AND_u1_u1_3897_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_3855_to_assign_stmt_3898/AND_u1_u1_3897_Update/$entry
      -- 	branch_block_stmt_2042/assign_stmt_3855_to_assign_stmt_3898/AND_u1_u1_3897_Update/cr
      -- 
    cp_elements(1178) <= cp_elements(1149);
    cr_15169_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1178), ack => AND_u1_u1_3897_inst_req_1); -- 
    -- CP-element group 1179 transition  input  bypass 
    -- predecessors 1177 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_3855_to_assign_stmt_3898/AND_u1_u1_3897_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3855_to_assign_stmt_3898/AND_u1_u1_3897_Sample/$exit
      -- 	branch_block_stmt_2042/assign_stmt_3855_to_assign_stmt_3898/AND_u1_u1_3897_Sample/ra
      -- 
    ra_15165_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => AND_u1_u1_3897_inst_ack_0, ack => cp_elements(1179)); -- 
    -- CP-element group 1180 transition  input  bypass 
    -- predecessors 1178 
    -- successors 1181 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_3855_to_assign_stmt_3898/AND_u1_u1_3897_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3855_to_assign_stmt_3898/AND_u1_u1_3897_Update/$exit
      -- 	branch_block_stmt_2042/assign_stmt_3855_to_assign_stmt_3898/AND_u1_u1_3897_Update/ca
      -- 
    ca_15170_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => AND_u1_u1_3897_inst_ack_1, ack => cp_elements(1180)); -- 
    -- CP-element group 1181 join  transition  bypass 
    -- predecessors 1157 1163 1180 
    -- successors 73 
    -- members (1) 
      -- 	branch_block_stmt_2042/assign_stmt_3855_to_assign_stmt_3898/$exit
      -- 
    cp_element_group_1181: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1181"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= cp_elements(1157) & cp_elements(1163) & cp_elements(1180);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1181), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1182 transition  place  dead  bypass 
    -- predecessors 73 
    -- successors 74 
    -- members (8) 
      -- 	branch_block_stmt_2042/if_stmt_3899__exit__
      -- 	branch_block_stmt_2042/merge_stmt_3905__entry__
      -- 	branch_block_stmt_2042/if_stmt_3899_dead_link/$entry
      -- 	branch_block_stmt_2042/if_stmt_3899_dead_link/$exit
      -- 	branch_block_stmt_2042/if_stmt_3899_dead_link/dead_transition
      -- 	branch_block_stmt_2042/merge_stmt_3905_dead_link/$entry
      -- 	branch_block_stmt_2042/merge_stmt_3905_dead_link/$exit
      -- 	branch_block_stmt_2042/merge_stmt_3905_dead_link/dead_transition
      -- 
    cp_elements(1182) <= false;
    -- CP-element group 1183 transition  output  bypass 
    -- predecessors 73 
    -- successors 1184 
    -- members (3) 
      -- 	branch_block_stmt_2042/if_stmt_3899_eval_test/$entry
      -- 	branch_block_stmt_2042/if_stmt_3899_eval_test/$exit
      -- 	branch_block_stmt_2042/if_stmt_3899_eval_test/branch_req
      -- 
    cp_elements(1183) <= cp_elements(73);
    branch_req_15178_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1183), ack => if_stmt_3899_branch_req_0); -- 
    -- CP-element group 1184 branch  place  bypass 
    -- predecessors 1183 
    -- successors 1185 1187 
    -- members (1) 
      -- 	branch_block_stmt_2042/R_orx_xcond11x_xi_3900_place
      -- 
    cp_elements(1184) <= cp_elements(1183);
    -- CP-element group 1185 transition  bypass 
    -- predecessors 1184 
    -- successors 1186 
    -- members (1) 
      -- 	branch_block_stmt_2042/if_stmt_3899_if_link/$entry
      -- 
    cp_elements(1185) <= cp_elements(1184);
    -- CP-element group 1186 transition  place  input  bypass 
    -- predecessors 1185 
    -- successors 74 
    -- members (9) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xpreheaderx_xi_udiv32x_xexitx_xix_xpreheader
      -- 	branch_block_stmt_2042/if_stmt_3899_if_link/$exit
      -- 	branch_block_stmt_2042/if_stmt_3899_if_link/if_choice_transition
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xpreheaderx_xi_udiv32x_xexitx_xix_xpreheader_PhiReq/$entry
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xpreheaderx_xi_udiv32x_xexitx_xix_xpreheader_PhiReq/$exit
      -- 	branch_block_stmt_2042/merge_stmt_3905_PhiReqMerge
      -- 	branch_block_stmt_2042/merge_stmt_3905_PhiAck/$entry
      -- 	branch_block_stmt_2042/merge_stmt_3905_PhiAck/$exit
      -- 	branch_block_stmt_2042/merge_stmt_3905_PhiAck/dummy
      -- 
    if_choice_transition_15183_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_3899_branch_ack_1, ack => cp_elements(1186)); -- 
    -- CP-element group 1187 transition  bypass 
    -- predecessors 1184 
    -- successors 1188 
    -- members (1) 
      -- 	branch_block_stmt_2042/if_stmt_3899_else_link/$entry
      -- 
    cp_elements(1187) <= cp_elements(1184);
    -- CP-element group 1188 transition  place  input  bypass 
    -- predecessors 1187 
    -- successors 2518 
    -- members (3) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xpreheaderx_xi_xx_xcritedgex_xi
      -- 	branch_block_stmt_2042/if_stmt_3899_else_link/$exit
      -- 	branch_block_stmt_2042/if_stmt_3899_else_link/else_choice_transition
      -- 
    else_choice_transition_15187_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_3899_branch_ack_0, ack => cp_elements(1188)); -- 
    -- CP-element group 1189 fork  transition  bypass 
    -- predecessors 75 
    -- successors 1190 1191 1194 1198 1201 1208 1211 1212 
    -- members (1) 
      -- 	branch_block_stmt_2042/assign_stmt_3927_to_assign_stmt_3958/$entry
      -- 
    cp_elements(1189) <= cp_elements(75);
    -- CP-element group 1190 transition  output  bypass 
    -- predecessors 1189 
    -- successors 1193 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_3927_to_assign_stmt_3958/SHL_u32_u32_3926_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_3927_to_assign_stmt_3958/SHL_u32_u32_3926_Update/$entry
      -- 	branch_block_stmt_2042/assign_stmt_3927_to_assign_stmt_3958/SHL_u32_u32_3926_Update/cr
      -- 
    cp_elements(1190) <= cp_elements(1189);
    cr_15209_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1190), ack => SHL_u32_u32_3926_inst_req_1); -- 
    -- CP-element group 1191 transition  output  bypass 
    -- predecessors 1189 
    -- successors 1192 
    -- members (7) 
      -- 	branch_block_stmt_2042/assign_stmt_3927_to_assign_stmt_3958/SHL_u32_u32_3926_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_3927_to_assign_stmt_3958/R_tempx_x012x_xi_3923_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_3927_to_assign_stmt_3958/R_tempx_x012x_xi_3923_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3927_to_assign_stmt_3958/R_tempx_x012x_xi_3923_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_3927_to_assign_stmt_3958/R_tempx_x012x_xi_3923_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3927_to_assign_stmt_3958/SHL_u32_u32_3926_Sample/$entry
      -- 	branch_block_stmt_2042/assign_stmt_3927_to_assign_stmt_3958/SHL_u32_u32_3926_Sample/rr
      -- 
    cp_elements(1191) <= cp_elements(1189);
    rr_15204_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1191), ack => SHL_u32_u32_3926_inst_req_0); -- 
    -- CP-element group 1192 transition  input  bypass 
    -- predecessors 1191 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_3927_to_assign_stmt_3958/SHL_u32_u32_3926_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3927_to_assign_stmt_3958/SHL_u32_u32_3926_Sample/$exit
      -- 	branch_block_stmt_2042/assign_stmt_3927_to_assign_stmt_3958/SHL_u32_u32_3926_Sample/ra
      -- 
    ra_15205_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => SHL_u32_u32_3926_inst_ack_0, ack => cp_elements(1192)); -- 
    -- CP-element group 1193 fork  transition  input  bypass 
    -- predecessors 1190 
    -- successors 1195 1202 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_3927_to_assign_stmt_3958/SHL_u32_u32_3926_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3927_to_assign_stmt_3958/SHL_u32_u32_3926_Update/$exit
      -- 	branch_block_stmt_2042/assign_stmt_3927_to_assign_stmt_3958/SHL_u32_u32_3926_Update/ca
      -- 
    ca_15210_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => SHL_u32_u32_3926_inst_ack_1, ack => cp_elements(1193)); -- 
    -- CP-element group 1194 transition  output  bypass 
    -- predecessors 1189 
    -- successors 1197 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_3927_to_assign_stmt_3958/AND_u32_u32_3932_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_3927_to_assign_stmt_3958/AND_u32_u32_3932_Update/$entry
      -- 	branch_block_stmt_2042/assign_stmt_3927_to_assign_stmt_3958/AND_u32_u32_3932_Update/cr
      -- 
    cp_elements(1194) <= cp_elements(1189);
    cr_15227_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1194), ack => AND_u32_u32_3932_inst_req_1); -- 
    -- CP-element group 1195 transition  output  bypass 
    -- predecessors 1193 
    -- successors 1196 
    -- members (7) 
      -- 	branch_block_stmt_2042/assign_stmt_3927_to_assign_stmt_3958/AND_u32_u32_3932_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_3927_to_assign_stmt_3958/R_iNsTr_256_3929_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_3927_to_assign_stmt_3958/R_iNsTr_256_3929_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3927_to_assign_stmt_3958/R_iNsTr_256_3929_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_3927_to_assign_stmt_3958/R_iNsTr_256_3929_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3927_to_assign_stmt_3958/AND_u32_u32_3932_Sample/$entry
      -- 	branch_block_stmt_2042/assign_stmt_3927_to_assign_stmt_3958/AND_u32_u32_3932_Sample/rr
      -- 
    cp_elements(1195) <= cp_elements(1193);
    rr_15222_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1195), ack => AND_u32_u32_3932_inst_req_0); -- 
    -- CP-element group 1196 transition  input  bypass 
    -- predecessors 1195 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_3927_to_assign_stmt_3958/AND_u32_u32_3932_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3927_to_assign_stmt_3958/AND_u32_u32_3932_Sample/$exit
      -- 	branch_block_stmt_2042/assign_stmt_3927_to_assign_stmt_3958/AND_u32_u32_3932_Sample/ra
      -- 
    ra_15223_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => AND_u32_u32_3932_inst_ack_0, ack => cp_elements(1196)); -- 
    -- CP-element group 1197 transition  input  output  bypass 
    -- predecessors 1194 
    -- successors 1199 
    -- members (10) 
      -- 	branch_block_stmt_2042/assign_stmt_3927_to_assign_stmt_3958/AND_u32_u32_3932_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3927_to_assign_stmt_3958/AND_u32_u32_3932_Update/$exit
      -- 	branch_block_stmt_2042/assign_stmt_3927_to_assign_stmt_3958/AND_u32_u32_3932_Update/ca
      -- 	branch_block_stmt_2042/assign_stmt_3927_to_assign_stmt_3958/EQ_u32_u1_3938_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_3927_to_assign_stmt_3958/R_iNsTr_257_3935_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_3927_to_assign_stmt_3958/R_iNsTr_257_3935_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3927_to_assign_stmt_3958/R_iNsTr_257_3935_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_3927_to_assign_stmt_3958/R_iNsTr_257_3935_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3927_to_assign_stmt_3958/EQ_u32_u1_3938_Sample/$entry
      -- 	branch_block_stmt_2042/assign_stmt_3927_to_assign_stmt_3958/EQ_u32_u1_3938_Sample/rr
      -- 
    ca_15228_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => AND_u32_u32_3932_inst_ack_1, ack => cp_elements(1197)); -- 
    rr_15240_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1197), ack => EQ_u32_u1_3938_inst_req_0); -- 
    -- CP-element group 1198 transition  output  bypass 
    -- predecessors 1189 
    -- successors 1200 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_3927_to_assign_stmt_3958/EQ_u32_u1_3938_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_3927_to_assign_stmt_3958/EQ_u32_u1_3938_Update/$entry
      -- 	branch_block_stmt_2042/assign_stmt_3927_to_assign_stmt_3958/EQ_u32_u1_3938_Update/cr
      -- 
    cp_elements(1198) <= cp_elements(1189);
    cr_15245_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1198), ack => EQ_u32_u1_3938_inst_req_1); -- 
    -- CP-element group 1199 transition  input  bypass 
    -- predecessors 1197 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_3927_to_assign_stmt_3958/EQ_u32_u1_3938_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3927_to_assign_stmt_3958/EQ_u32_u1_3938_Sample/$exit
      -- 	branch_block_stmt_2042/assign_stmt_3927_to_assign_stmt_3958/EQ_u32_u1_3938_Sample/ra
      -- 
    ra_15241_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u32_u1_3938_inst_ack_0, ack => cp_elements(1199)); -- 
    -- CP-element group 1200 transition  input  bypass 
    -- predecessors 1198 
    -- successors 1207 
    -- members (7) 
      -- 	branch_block_stmt_2042/assign_stmt_3927_to_assign_stmt_3958/EQ_u32_u1_3938_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3927_to_assign_stmt_3958/EQ_u32_u1_3938_Update/$exit
      -- 	branch_block_stmt_2042/assign_stmt_3927_to_assign_stmt_3958/EQ_u32_u1_3938_Update/ca
      -- 	branch_block_stmt_2042/assign_stmt_3927_to_assign_stmt_3958/R_iNsTr_258_3949_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_3927_to_assign_stmt_3958/R_iNsTr_258_3949_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3927_to_assign_stmt_3958/R_iNsTr_258_3949_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_3927_to_assign_stmt_3958/R_iNsTr_258_3949_update_completed_
      -- 
    ca_15246_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u32_u1_3938_inst_ack_1, ack => cp_elements(1200)); -- 
    -- CP-element group 1201 transition  output  bypass 
    -- predecessors 1189 
    -- successors 1206 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_3927_to_assign_stmt_3958/NEQ_i32_u1_3946_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_3927_to_assign_stmt_3958/NEQ_i32_u1_3946_Update/$entry
      -- 	branch_block_stmt_2042/assign_stmt_3927_to_assign_stmt_3958/NEQ_i32_u1_3946_Update/cr
      -- 
    cp_elements(1201) <= cp_elements(1189);
    cr_15277_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1201), ack => NEQ_i32_u1_3946_inst_req_1); -- 
    -- CP-element group 1202 transition  output  bypass 
    -- predecessors 1193 
    -- successors 1203 
    -- members (7) 
      -- 	branch_block_stmt_2042/assign_stmt_3927_to_assign_stmt_3958/type_cast_3942_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_3927_to_assign_stmt_3958/R_iNsTr_256_3941_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_3927_to_assign_stmt_3958/R_iNsTr_256_3941_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3927_to_assign_stmt_3958/R_iNsTr_256_3941_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_3927_to_assign_stmt_3958/R_iNsTr_256_3941_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3927_to_assign_stmt_3958/type_cast_3942_Sample/$entry
      -- 	branch_block_stmt_2042/assign_stmt_3927_to_assign_stmt_3958/type_cast_3942_Sample/rr
      -- 
    cp_elements(1202) <= cp_elements(1193);
    rr_15262_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1202), ack => type_cast_3942_inst_req_0); -- 
    -- CP-element group 1203 transition  input  output  bypass 
    -- predecessors 1202 
    -- successors 1204 
    -- members (6) 
      -- 	branch_block_stmt_2042/assign_stmt_3927_to_assign_stmt_3958/type_cast_3942_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3927_to_assign_stmt_3958/type_cast_3942_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_3927_to_assign_stmt_3958/type_cast_3942_Sample/$exit
      -- 	branch_block_stmt_2042/assign_stmt_3927_to_assign_stmt_3958/type_cast_3942_Sample/ra
      -- 	branch_block_stmt_2042/assign_stmt_3927_to_assign_stmt_3958/type_cast_3942_Update/$entry
      -- 	branch_block_stmt_2042/assign_stmt_3927_to_assign_stmt_3958/type_cast_3942_Update/cr
      -- 
    ra_15263_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3942_inst_ack_0, ack => cp_elements(1203)); -- 
    cr_15267_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1203), ack => type_cast_3942_inst_req_1); -- 
    -- CP-element group 1204 transition  input  output  bypass 
    -- predecessors 1203 
    -- successors 1205 
    -- members (6) 
      -- 	branch_block_stmt_2042/assign_stmt_3927_to_assign_stmt_3958/NEQ_i32_u1_3946_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_3927_to_assign_stmt_3958/type_cast_3942_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3927_to_assign_stmt_3958/type_cast_3942_Update/$exit
      -- 	branch_block_stmt_2042/assign_stmt_3927_to_assign_stmt_3958/type_cast_3942_Update/ca
      -- 	branch_block_stmt_2042/assign_stmt_3927_to_assign_stmt_3958/NEQ_i32_u1_3946_Sample/$entry
      -- 	branch_block_stmt_2042/assign_stmt_3927_to_assign_stmt_3958/NEQ_i32_u1_3946_Sample/rr
      -- 
    ca_15268_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3942_inst_ack_1, ack => cp_elements(1204)); -- 
    rr_15272_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1204), ack => NEQ_i32_u1_3946_inst_req_0); -- 
    -- CP-element group 1205 transition  input  bypass 
    -- predecessors 1204 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_3927_to_assign_stmt_3958/NEQ_i32_u1_3946_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3927_to_assign_stmt_3958/NEQ_i32_u1_3946_Sample/$exit
      -- 	branch_block_stmt_2042/assign_stmt_3927_to_assign_stmt_3958/NEQ_i32_u1_3946_Sample/ra
      -- 
    ra_15273_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => NEQ_i32_u1_3946_inst_ack_0, ack => cp_elements(1205)); -- 
    -- CP-element group 1206 transition  input  bypass 
    -- predecessors 1201 
    -- successors 1207 
    -- members (7) 
      -- 	branch_block_stmt_2042/assign_stmt_3927_to_assign_stmt_3958/NEQ_i32_u1_3946_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3927_to_assign_stmt_3958/NEQ_i32_u1_3946_Update/$exit
      -- 	branch_block_stmt_2042/assign_stmt_3927_to_assign_stmt_3958/NEQ_i32_u1_3946_Update/ca
      -- 	branch_block_stmt_2042/assign_stmt_3927_to_assign_stmt_3958/R_iNsTr_259_3950_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_3927_to_assign_stmt_3958/R_iNsTr_259_3950_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3927_to_assign_stmt_3958/R_iNsTr_259_3950_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_3927_to_assign_stmt_3958/R_iNsTr_259_3950_update_completed_
      -- 
    ca_15278_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => NEQ_i32_u1_3946_inst_ack_1, ack => cp_elements(1206)); -- 
    -- CP-element group 1207 join  transition  output  bypass 
    -- predecessors 1200 1206 
    -- successors 1209 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_3927_to_assign_stmt_3958/AND_u1_u1_3951_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_3927_to_assign_stmt_3958/AND_u1_u1_3951_Sample/$entry
      -- 	branch_block_stmt_2042/assign_stmt_3927_to_assign_stmt_3958/AND_u1_u1_3951_Sample/rr
      -- 
    cp_element_group_1207: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1207"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1200) & cp_elements(1206);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1207), clk => clk, reset => reset); --
    end block;
    rr_15294_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1207), ack => AND_u1_u1_3951_inst_req_0); -- 
    -- CP-element group 1208 transition  output  bypass 
    -- predecessors 1189 
    -- successors 1210 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_3927_to_assign_stmt_3958/AND_u1_u1_3951_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_3927_to_assign_stmt_3958/AND_u1_u1_3951_Update/$entry
      -- 	branch_block_stmt_2042/assign_stmt_3927_to_assign_stmt_3958/AND_u1_u1_3951_Update/cr
      -- 
    cp_elements(1208) <= cp_elements(1189);
    cr_15299_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1208), ack => AND_u1_u1_3951_inst_req_1); -- 
    -- CP-element group 1209 transition  input  bypass 
    -- predecessors 1207 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_3927_to_assign_stmt_3958/AND_u1_u1_3951_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3927_to_assign_stmt_3958/AND_u1_u1_3951_Sample/$exit
      -- 	branch_block_stmt_2042/assign_stmt_3927_to_assign_stmt_3958/AND_u1_u1_3951_Sample/ra
      -- 
    ra_15295_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => AND_u1_u1_3951_inst_ack_0, ack => cp_elements(1209)); -- 
    -- CP-element group 1210 transition  input  bypass 
    -- predecessors 1208 
    -- successors 1215 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_3927_to_assign_stmt_3958/AND_u1_u1_3951_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3927_to_assign_stmt_3958/AND_u1_u1_3951_Update/$exit
      -- 	branch_block_stmt_2042/assign_stmt_3927_to_assign_stmt_3958/AND_u1_u1_3951_Update/ca
      -- 
    ca_15300_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => AND_u1_u1_3951_inst_ack_1, ack => cp_elements(1210)); -- 
    -- CP-element group 1211 transition  output  bypass 
    -- predecessors 1189 
    -- successors 1214 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_3927_to_assign_stmt_3958/ADD_u32_u32_3957_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_3927_to_assign_stmt_3958/ADD_u32_u32_3957_Update/$entry
      -- 	branch_block_stmt_2042/assign_stmt_3927_to_assign_stmt_3958/ADD_u32_u32_3957_Update/cr
      -- 
    cp_elements(1211) <= cp_elements(1189);
    cr_15317_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1211), ack => ADD_u32_u32_3957_inst_req_1); -- 
    -- CP-element group 1212 transition  output  bypass 
    -- predecessors 1189 
    -- successors 1213 
    -- members (7) 
      -- 	branch_block_stmt_2042/assign_stmt_3927_to_assign_stmt_3958/ADD_u32_u32_3957_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_3927_to_assign_stmt_3958/R_iNsTr_255_3954_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_3927_to_assign_stmt_3958/R_iNsTr_255_3954_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3927_to_assign_stmt_3958/R_iNsTr_255_3954_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_3927_to_assign_stmt_3958/R_iNsTr_255_3954_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3927_to_assign_stmt_3958/ADD_u32_u32_3957_Sample/$entry
      -- 	branch_block_stmt_2042/assign_stmt_3927_to_assign_stmt_3958/ADD_u32_u32_3957_Sample/rr
      -- 
    cp_elements(1212) <= cp_elements(1189);
    rr_15312_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1212), ack => ADD_u32_u32_3957_inst_req_0); -- 
    -- CP-element group 1213 transition  input  bypass 
    -- predecessors 1212 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_3927_to_assign_stmt_3958/ADD_u32_u32_3957_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3927_to_assign_stmt_3958/ADD_u32_u32_3957_Sample/$exit
      -- 	branch_block_stmt_2042/assign_stmt_3927_to_assign_stmt_3958/ADD_u32_u32_3957_Sample/ra
      -- 
    ra_15313_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u32_u32_3957_inst_ack_0, ack => cp_elements(1213)); -- 
    -- CP-element group 1214 transition  input  bypass 
    -- predecessors 1211 
    -- successors 1215 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_3927_to_assign_stmt_3958/ADD_u32_u32_3957_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3927_to_assign_stmt_3958/ADD_u32_u32_3957_Update/$exit
      -- 	branch_block_stmt_2042/assign_stmt_3927_to_assign_stmt_3958/ADD_u32_u32_3957_Update/ca
      -- 
    ca_15318_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u32_u32_3957_inst_ack_1, ack => cp_elements(1214)); -- 
    -- CP-element group 1215 join  transition  bypass 
    -- predecessors 1210 1214 
    -- successors 76 
    -- members (1) 
      -- 	branch_block_stmt_2042/assign_stmt_3927_to_assign_stmt_3958/$exit
      -- 
    cp_element_group_1215: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1215"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1210) & cp_elements(1214);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1215), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1216 transition  place  dead  bypass 
    -- predecessors 76 
    -- successors 77 
    -- members (8) 
      -- 	branch_block_stmt_2042/if_stmt_3959__exit__
      -- 	branch_block_stmt_2042/merge_stmt_3965__entry__
      -- 	branch_block_stmt_2042/if_stmt_3959_dead_link/$entry
      -- 	branch_block_stmt_2042/if_stmt_3959_dead_link/$exit
      -- 	branch_block_stmt_2042/if_stmt_3959_dead_link/dead_transition
      -- 	branch_block_stmt_2042/merge_stmt_3965_dead_link/$entry
      -- 	branch_block_stmt_2042/merge_stmt_3965_dead_link/$exit
      -- 	branch_block_stmt_2042/merge_stmt_3965_dead_link/dead_transition
      -- 
    cp_elements(1216) <= false;
    -- CP-element group 1217 transition  output  bypass 
    -- predecessors 76 
    -- successors 1218 
    -- members (3) 
      -- 	branch_block_stmt_2042/if_stmt_3959_eval_test/$entry
      -- 	branch_block_stmt_2042/if_stmt_3959_eval_test/$exit
      -- 	branch_block_stmt_2042/if_stmt_3959_eval_test/branch_req
      -- 
    cp_elements(1217) <= cp_elements(76);
    branch_req_15326_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1217), ack => if_stmt_3959_branch_req_0); -- 
    -- CP-element group 1218 branch  place  bypass 
    -- predecessors 1217 
    -- successors 1219 1221 
    -- members (1) 
      -- 	branch_block_stmt_2042/R_orx_xcondx_xi_3960_place
      -- 
    cp_elements(1218) <= cp_elements(1217);
    -- CP-element group 1219 transition  bypass 
    -- predecessors 1218 
    -- successors 1220 
    -- members (1) 
      -- 	branch_block_stmt_2042/if_stmt_3959_if_link/$entry
      -- 
    cp_elements(1219) <= cp_elements(1218);
    -- CP-element group 1220 transition  place  input  bypass 
    -- predecessors 1219 
    -- successors 2456 
    -- members (3) 
      -- 	branch_block_stmt_2042/if_stmt_3959_if_link/$exit
      -- 	branch_block_stmt_2042/if_stmt_3959_if_link/if_choice_transition
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xi_udiv32x_xexitx_xi
      -- 
    if_choice_transition_15331_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_3959_branch_ack_1, ack => cp_elements(1220)); -- 
    -- CP-element group 1221 transition  bypass 
    -- predecessors 1218 
    -- successors 1222 
    -- members (1) 
      -- 	branch_block_stmt_2042/if_stmt_3959_else_link/$entry
      -- 
    cp_elements(1221) <= cp_elements(1218);
    -- CP-element group 1222 transition  place  input  bypass 
    -- predecessors 1221 
    -- successors 2499 
    -- members (3) 
      -- 	branch_block_stmt_2042/if_stmt_3959_else_link/$exit
      -- 	branch_block_stmt_2042/if_stmt_3959_else_link/else_choice_transition
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xi_udiv32x_xexitx_xx_xcritedge_crit_edgex_xi
      -- 
    else_choice_transition_15335_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_3959_branch_ack_0, ack => cp_elements(1222)); -- 
    -- CP-element group 1223 fork  transition  bypass 
    -- predecessors 77 
    -- successors 1224 1225 1229 1230 
    -- members (1) 
      -- 	branch_block_stmt_2042/assign_stmt_3980_to_assign_stmt_3985/$entry
      -- 
    cp_elements(1223) <= cp_elements(77);
    -- CP-element group 1224 transition  output  bypass 
    -- predecessors 1223 
    -- successors 1227 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_3980_to_assign_stmt_3985/ADD_u32_u32_3979_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_3980_to_assign_stmt_3985/ADD_u32_u32_3979_Update/$entry
      -- 	branch_block_stmt_2042/assign_stmt_3980_to_assign_stmt_3985/ADD_u32_u32_3979_Update/cr
      -- 
    cp_elements(1224) <= cp_elements(1223);
    cr_15357_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1224), ack => ADD_u32_u32_3979_inst_req_1); -- 
    -- CP-element group 1225 transition  output  bypass 
    -- predecessors 1223 
    -- successors 1226 
    -- members (7) 
      -- 	branch_block_stmt_2042/assign_stmt_3980_to_assign_stmt_3985/ADD_u32_u32_3979_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_3980_to_assign_stmt_3985/R_iNsTr_240_3976_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_3980_to_assign_stmt_3985/R_iNsTr_240_3976_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3980_to_assign_stmt_3985/R_iNsTr_240_3976_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_3980_to_assign_stmt_3985/R_iNsTr_240_3976_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3980_to_assign_stmt_3985/ADD_u32_u32_3979_Sample/$entry
      -- 	branch_block_stmt_2042/assign_stmt_3980_to_assign_stmt_3985/ADD_u32_u32_3979_Sample/rr
      -- 
    cp_elements(1225) <= cp_elements(1223);
    rr_15352_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1225), ack => ADD_u32_u32_3979_inst_req_0); -- 
    -- CP-element group 1226 transition  input  bypass 
    -- predecessors 1225 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_3980_to_assign_stmt_3985/ADD_u32_u32_3979_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3980_to_assign_stmt_3985/ADD_u32_u32_3979_Sample/$exit
      -- 	branch_block_stmt_2042/assign_stmt_3980_to_assign_stmt_3985/ADD_u32_u32_3979_Sample/ra
      -- 
    ra_15353_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u32_u32_3979_inst_ack_0, ack => cp_elements(1226)); -- 
    -- CP-element group 1227 transition  input  bypass 
    -- predecessors 1224 
    -- successors 1228 
    -- members (7) 
      -- 	branch_block_stmt_2042/assign_stmt_3980_to_assign_stmt_3985/ADD_u32_u32_3979_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3980_to_assign_stmt_3985/ADD_u32_u32_3979_Update/$exit
      -- 	branch_block_stmt_2042/assign_stmt_3980_to_assign_stmt_3985/ADD_u32_u32_3979_Update/ca
      -- 	branch_block_stmt_2042/assign_stmt_3980_to_assign_stmt_3985/R_tmp25x_xi_3982_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_3980_to_assign_stmt_3985/R_tmp25x_xi_3982_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3980_to_assign_stmt_3985/R_tmp25x_xi_3982_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_3980_to_assign_stmt_3985/R_tmp25x_xi_3982_update_completed_
      -- 
    ca_15358_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u32_u32_3979_inst_ack_1, ack => cp_elements(1227)); -- 
    -- CP-element group 1228 join  transition  output  bypass 
    -- predecessors 1227 1230 
    -- successors 1231 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_3980_to_assign_stmt_3985/SUB_u32_u32_3984_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_3980_to_assign_stmt_3985/SUB_u32_u32_3984_Sample/$entry
      -- 	branch_block_stmt_2042/assign_stmt_3980_to_assign_stmt_3985/SUB_u32_u32_3984_Sample/rr
      -- 
    cp_element_group_1228: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1228"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1227) & cp_elements(1230);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1228), clk => clk, reset => reset); --
    end block;
    rr_15374_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1228), ack => SUB_u32_u32_3984_inst_req_0); -- 
    -- CP-element group 1229 transition  output  bypass 
    -- predecessors 1223 
    -- successors 1232 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_3980_to_assign_stmt_3985/SUB_u32_u32_3984_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_3980_to_assign_stmt_3985/SUB_u32_u32_3984_Update/$entry
      -- 	branch_block_stmt_2042/assign_stmt_3980_to_assign_stmt_3985/SUB_u32_u32_3984_Update/cr
      -- 
    cp_elements(1229) <= cp_elements(1223);
    cr_15379_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1229), ack => SUB_u32_u32_3984_inst_req_1); -- 
    -- CP-element group 1230 transition  bypass 
    -- predecessors 1223 
    -- successors 1228 
    -- members (4) 
      -- 	branch_block_stmt_2042/assign_stmt_3980_to_assign_stmt_3985/R_xx_xlcssa_3983_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_3980_to_assign_stmt_3985/R_xx_xlcssa_3983_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3980_to_assign_stmt_3985/R_xx_xlcssa_3983_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_3980_to_assign_stmt_3985/R_xx_xlcssa_3983_update_completed_
      -- 
    cp_elements(1230) <= cp_elements(1223);
    -- CP-element group 1231 transition  input  bypass 
    -- predecessors 1228 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_3980_to_assign_stmt_3985/SUB_u32_u32_3984_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3980_to_assign_stmt_3985/SUB_u32_u32_3984_Sample/$exit
      -- 	branch_block_stmt_2042/assign_stmt_3980_to_assign_stmt_3985/SUB_u32_u32_3984_Sample/ra
      -- 
    ra_15375_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => SUB_u32_u32_3984_inst_ack_0, ack => cp_elements(1231)); -- 
    -- CP-element group 1232 transition  place  input  bypass 
    -- predecessors 1229 
    -- successors 2544 
    -- members (6) 
      -- 	branch_block_stmt_2042/assign_stmt_3980_to_assign_stmt_3985__exit__
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xx_xcritedge_crit_edgex_xi_xx_xcritedgex_xi
      -- 	branch_block_stmt_2042/assign_stmt_3980_to_assign_stmt_3985/$exit
      -- 	branch_block_stmt_2042/assign_stmt_3980_to_assign_stmt_3985/SUB_u32_u32_3984_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_3980_to_assign_stmt_3985/SUB_u32_u32_3984_Update/$exit
      -- 	branch_block_stmt_2042/assign_stmt_3980_to_assign_stmt_3985/SUB_u32_u32_3984_Update/ca
      -- 
    ca_15380_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => SUB_u32_u32_3984_inst_ack_1, ack => cp_elements(1232)); -- 
    -- CP-element group 1233 fork  transition  bypass 
    -- predecessors 78 
    -- successors 1234 1235 1238 1239 1242 1246 1247 1251 1254 
    -- members (1) 
      -- 	branch_block_stmt_2042/assign_stmt_4006_to_assign_stmt_4032/$entry
      -- 
    cp_elements(1233) <= cp_elements(78);
    -- CP-element group 1234 transition  output  bypass 
    -- predecessors 1233 
    -- successors 1237 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_4006_to_assign_stmt_4032/AND_u32_u32_4005_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_4006_to_assign_stmt_4032/AND_u32_u32_4005_Update/$entry
      -- 	branch_block_stmt_2042/assign_stmt_4006_to_assign_stmt_4032/AND_u32_u32_4005_Update/cr
      -- 
    cp_elements(1234) <= cp_elements(1233);
    cr_15400_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1234), ack => AND_u32_u32_4005_inst_req_1); -- 
    -- CP-element group 1235 transition  output  bypass 
    -- predecessors 1233 
    -- successors 1236 
    -- members (7) 
      -- 	branch_block_stmt_2042/assign_stmt_4006_to_assign_stmt_4032/AND_u32_u32_4005_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_4006_to_assign_stmt_4032/R_tempx_x0x_xlcssax_xi_4002_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_4006_to_assign_stmt_4032/R_tempx_x0x_xlcssax_xi_4002_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_4006_to_assign_stmt_4032/R_tempx_x0x_xlcssax_xi_4002_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_4006_to_assign_stmt_4032/R_tempx_x0x_xlcssax_xi_4002_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_4006_to_assign_stmt_4032/AND_u32_u32_4005_Sample/$entry
      -- 	branch_block_stmt_2042/assign_stmt_4006_to_assign_stmt_4032/AND_u32_u32_4005_Sample/rr
      -- 
    cp_elements(1235) <= cp_elements(1233);
    rr_15395_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1235), ack => AND_u32_u32_4005_inst_req_0); -- 
    -- CP-element group 1236 transition  input  bypass 
    -- predecessors 1235 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_4006_to_assign_stmt_4032/AND_u32_u32_4005_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_4006_to_assign_stmt_4032/AND_u32_u32_4005_Sample/$exit
      -- 	branch_block_stmt_2042/assign_stmt_4006_to_assign_stmt_4032/AND_u32_u32_4005_Sample/ra
      -- 
    ra_15396_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => AND_u32_u32_4005_inst_ack_0, ack => cp_elements(1236)); -- 
    -- CP-element group 1237 transition  input  bypass 
    -- predecessors 1234 
    -- successors 1250 
    -- members (7) 
      -- 	branch_block_stmt_2042/assign_stmt_4006_to_assign_stmt_4032/AND_u32_u32_4005_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_4006_to_assign_stmt_4032/AND_u32_u32_4005_Update/$exit
      -- 	branch_block_stmt_2042/assign_stmt_4006_to_assign_stmt_4032/AND_u32_u32_4005_Update/ca
      -- 	branch_block_stmt_2042/assign_stmt_4006_to_assign_stmt_4032/R_iNsTr_249_4026_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_4006_to_assign_stmt_4032/R_iNsTr_249_4026_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_4006_to_assign_stmt_4032/R_iNsTr_249_4026_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_4006_to_assign_stmt_4032/R_iNsTr_249_4026_update_completed_
      -- 
    ca_15401_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => AND_u32_u32_4005_inst_ack_1, ack => cp_elements(1237)); -- 
    -- CP-element group 1238 transition  output  bypass 
    -- predecessors 1233 
    -- successors 1241 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_4006_to_assign_stmt_4032/SHL_u32_u32_4011_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_4006_to_assign_stmt_4032/SHL_u32_u32_4011_Update/$entry
      -- 	branch_block_stmt_2042/assign_stmt_4006_to_assign_stmt_4032/SHL_u32_u32_4011_Update/cr
      -- 
    cp_elements(1238) <= cp_elements(1233);
    cr_15418_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1238), ack => SHL_u32_u32_4011_inst_req_1); -- 
    -- CP-element group 1239 transition  output  bypass 
    -- predecessors 1233 
    -- successors 1240 
    -- members (7) 
      -- 	branch_block_stmt_2042/assign_stmt_4006_to_assign_stmt_4032/SHL_u32_u32_4011_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_4006_to_assign_stmt_4032/R_expx_x0x_xlcssax_xi_4008_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_4006_to_assign_stmt_4032/R_expx_x0x_xlcssax_xi_4008_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_4006_to_assign_stmt_4032/R_expx_x0x_xlcssax_xi_4008_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_4006_to_assign_stmt_4032/R_expx_x0x_xlcssax_xi_4008_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_4006_to_assign_stmt_4032/SHL_u32_u32_4011_Sample/$entry
      -- 	branch_block_stmt_2042/assign_stmt_4006_to_assign_stmt_4032/SHL_u32_u32_4011_Sample/rr
      -- 
    cp_elements(1239) <= cp_elements(1233);
    rr_15413_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1239), ack => SHL_u32_u32_4011_inst_req_0); -- 
    -- CP-element group 1240 transition  input  bypass 
    -- predecessors 1239 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_4006_to_assign_stmt_4032/SHL_u32_u32_4011_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_4006_to_assign_stmt_4032/SHL_u32_u32_4011_Sample/$exit
      -- 	branch_block_stmt_2042/assign_stmt_4006_to_assign_stmt_4032/SHL_u32_u32_4011_Sample/ra
      -- 
    ra_15414_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => SHL_u32_u32_4011_inst_ack_0, ack => cp_elements(1240)); -- 
    -- CP-element group 1241 transition  input  output  bypass 
    -- predecessors 1238 
    -- successors 1243 
    -- members (10) 
      -- 	branch_block_stmt_2042/assign_stmt_4006_to_assign_stmt_4032/SHL_u32_u32_4011_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_4006_to_assign_stmt_4032/SHL_u32_u32_4011_Update/$exit
      -- 	branch_block_stmt_2042/assign_stmt_4006_to_assign_stmt_4032/SHL_u32_u32_4011_Update/ca
      -- 	branch_block_stmt_2042/assign_stmt_4006_to_assign_stmt_4032/ADD_u32_u32_4017_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_4006_to_assign_stmt_4032/R_iNsTr_250_4014_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_4006_to_assign_stmt_4032/R_iNsTr_250_4014_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_4006_to_assign_stmt_4032/R_iNsTr_250_4014_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_4006_to_assign_stmt_4032/R_iNsTr_250_4014_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_4006_to_assign_stmt_4032/ADD_u32_u32_4017_Sample/$entry
      -- 	branch_block_stmt_2042/assign_stmt_4006_to_assign_stmt_4032/ADD_u32_u32_4017_Sample/rr
      -- 
    ca_15419_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => SHL_u32_u32_4011_inst_ack_1, ack => cp_elements(1241)); -- 
    rr_15431_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1241), ack => ADD_u32_u32_4017_inst_req_0); -- 
    -- CP-element group 1242 transition  output  bypass 
    -- predecessors 1233 
    -- successors 1244 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_4006_to_assign_stmt_4032/ADD_u32_u32_4017_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_4006_to_assign_stmt_4032/ADD_u32_u32_4017_Update/$entry
      -- 	branch_block_stmt_2042/assign_stmt_4006_to_assign_stmt_4032/ADD_u32_u32_4017_Update/cr
      -- 
    cp_elements(1242) <= cp_elements(1233);
    cr_15436_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1242), ack => ADD_u32_u32_4017_inst_req_1); -- 
    -- CP-element group 1243 transition  input  bypass 
    -- predecessors 1241 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_4006_to_assign_stmt_4032/ADD_u32_u32_4017_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_4006_to_assign_stmt_4032/ADD_u32_u32_4017_Sample/$exit
      -- 	branch_block_stmt_2042/assign_stmt_4006_to_assign_stmt_4032/ADD_u32_u32_4017_Sample/ra
      -- 
    ra_15432_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u32_u32_4017_inst_ack_0, ack => cp_elements(1243)); -- 
    -- CP-element group 1244 transition  input  bypass 
    -- predecessors 1242 
    -- successors 1245 
    -- members (7) 
      -- 	branch_block_stmt_2042/assign_stmt_4006_to_assign_stmt_4032/ADD_u32_u32_4017_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_4006_to_assign_stmt_4032/ADD_u32_u32_4017_Update/$exit
      -- 	branch_block_stmt_2042/assign_stmt_4006_to_assign_stmt_4032/ADD_u32_u32_4017_Update/ca
      -- 	branch_block_stmt_2042/assign_stmt_4006_to_assign_stmt_4032/R_iNsTr_251_4020_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_4006_to_assign_stmt_4032/R_iNsTr_251_4020_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_4006_to_assign_stmt_4032/R_iNsTr_251_4020_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_4006_to_assign_stmt_4032/R_iNsTr_251_4020_update_completed_
      -- 
    ca_15437_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u32_u32_4017_inst_ack_1, ack => cp_elements(1244)); -- 
    -- CP-element group 1245 join  transition  output  bypass 
    -- predecessors 1244 1247 
    -- successors 1248 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_4006_to_assign_stmt_4032/OR_u32_u32_4022_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_4006_to_assign_stmt_4032/OR_u32_u32_4022_Sample/$entry
      -- 	branch_block_stmt_2042/assign_stmt_4006_to_assign_stmt_4032/OR_u32_u32_4022_Sample/rr
      -- 
    cp_element_group_1245: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1245"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1244) & cp_elements(1247);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1245), clk => clk, reset => reset); --
    end block;
    rr_15453_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1245), ack => OR_u32_u32_4022_inst_req_0); -- 
    -- CP-element group 1246 transition  output  bypass 
    -- predecessors 1233 
    -- successors 1249 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_4006_to_assign_stmt_4032/OR_u32_u32_4022_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_4006_to_assign_stmt_4032/OR_u32_u32_4022_Update/$entry
      -- 	branch_block_stmt_2042/assign_stmt_4006_to_assign_stmt_4032/OR_u32_u32_4022_Update/cr
      -- 
    cp_elements(1246) <= cp_elements(1233);
    cr_15458_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1246), ack => OR_u32_u32_4022_inst_req_1); -- 
    -- CP-element group 1247 transition  bypass 
    -- predecessors 1233 
    -- successors 1245 
    -- members (4) 
      -- 	branch_block_stmt_2042/assign_stmt_4006_to_assign_stmt_4032/R_iNsTr_239_4021_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_4006_to_assign_stmt_4032/R_iNsTr_239_4021_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_4006_to_assign_stmt_4032/R_iNsTr_239_4021_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_4006_to_assign_stmt_4032/R_iNsTr_239_4021_update_completed_
      -- 
    cp_elements(1247) <= cp_elements(1233);
    -- CP-element group 1248 transition  input  bypass 
    -- predecessors 1245 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_4006_to_assign_stmt_4032/OR_u32_u32_4022_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_4006_to_assign_stmt_4032/OR_u32_u32_4022_Sample/$exit
      -- 	branch_block_stmt_2042/assign_stmt_4006_to_assign_stmt_4032/OR_u32_u32_4022_Sample/ra
      -- 
    ra_15454_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => OR_u32_u32_4022_inst_ack_0, ack => cp_elements(1248)); -- 
    -- CP-element group 1249 transition  input  bypass 
    -- predecessors 1246 
    -- successors 1250 
    -- members (7) 
      -- 	branch_block_stmt_2042/assign_stmt_4006_to_assign_stmt_4032/OR_u32_u32_4022_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_4006_to_assign_stmt_4032/OR_u32_u32_4022_Update/$exit
      -- 	branch_block_stmt_2042/assign_stmt_4006_to_assign_stmt_4032/OR_u32_u32_4022_Update/ca
      -- 	branch_block_stmt_2042/assign_stmt_4006_to_assign_stmt_4032/R_iNsTr_252_4025_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_4006_to_assign_stmt_4032/R_iNsTr_252_4025_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_4006_to_assign_stmt_4032/R_iNsTr_252_4025_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_4006_to_assign_stmt_4032/R_iNsTr_252_4025_update_completed_
      -- 
    ca_15459_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => OR_u32_u32_4022_inst_ack_1, ack => cp_elements(1249)); -- 
    -- CP-element group 1250 join  transition  output  bypass 
    -- predecessors 1237 1249 
    -- successors 1252 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_4006_to_assign_stmt_4032/OR_u32_u32_4027_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_4006_to_assign_stmt_4032/OR_u32_u32_4027_Sample/$entry
      -- 	branch_block_stmt_2042/assign_stmt_4006_to_assign_stmt_4032/OR_u32_u32_4027_Sample/rr
      -- 
    cp_element_group_1250: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1250"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1237) & cp_elements(1249);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1250), clk => clk, reset => reset); --
    end block;
    rr_15475_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1250), ack => OR_u32_u32_4027_inst_req_0); -- 
    -- CP-element group 1251 transition  output  bypass 
    -- predecessors 1233 
    -- successors 1253 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_4006_to_assign_stmt_4032/OR_u32_u32_4027_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_4006_to_assign_stmt_4032/OR_u32_u32_4027_Update/$entry
      -- 	branch_block_stmt_2042/assign_stmt_4006_to_assign_stmt_4032/OR_u32_u32_4027_Update/cr
      -- 
    cp_elements(1251) <= cp_elements(1233);
    cr_15480_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1251), ack => OR_u32_u32_4027_inst_req_1); -- 
    -- CP-element group 1252 transition  input  bypass 
    -- predecessors 1250 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_4006_to_assign_stmt_4032/OR_u32_u32_4027_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_4006_to_assign_stmt_4032/OR_u32_u32_4027_Sample/$exit
      -- 	branch_block_stmt_2042/assign_stmt_4006_to_assign_stmt_4032/OR_u32_u32_4027_Sample/ra
      -- 
    ra_15476_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => OR_u32_u32_4027_inst_ack_0, ack => cp_elements(1252)); -- 
    -- CP-element group 1253 transition  input  output  bypass 
    -- predecessors 1251 
    -- successors 1255 
    -- members (10) 
      -- 	branch_block_stmt_2042/assign_stmt_4006_to_assign_stmt_4032/type_cast_4031_Sample/rr
      -- 	branch_block_stmt_2042/assign_stmt_4006_to_assign_stmt_4032/type_cast_4031_Sample/$entry
      -- 	branch_block_stmt_2042/assign_stmt_4006_to_assign_stmt_4032/R_iNsTr_253_4030_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_4006_to_assign_stmt_4032/OR_u32_u32_4027_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_4006_to_assign_stmt_4032/OR_u32_u32_4027_Update/$exit
      -- 	branch_block_stmt_2042/assign_stmt_4006_to_assign_stmt_4032/OR_u32_u32_4027_Update/ca
      -- 	branch_block_stmt_2042/assign_stmt_4006_to_assign_stmt_4032/type_cast_4031_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_4006_to_assign_stmt_4032/R_iNsTr_253_4030_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_4006_to_assign_stmt_4032/R_iNsTr_253_4030_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_4006_to_assign_stmt_4032/R_iNsTr_253_4030_update_start_
      -- 
    ca_15481_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => OR_u32_u32_4027_inst_ack_1, ack => cp_elements(1253)); -- 
    rr_15493_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1253), ack => type_cast_4031_inst_req_0); -- 
    -- CP-element group 1254 transition  output  bypass 
    -- predecessors 1233 
    -- successors 1256 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_4006_to_assign_stmt_4032/type_cast_4031_Update/cr
      -- 	branch_block_stmt_2042/assign_stmt_4006_to_assign_stmt_4032/type_cast_4031_Update/$entry
      -- 	branch_block_stmt_2042/assign_stmt_4006_to_assign_stmt_4032/type_cast_4031_update_start_
      -- 
    cp_elements(1254) <= cp_elements(1233);
    cr_15498_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1254), ack => type_cast_4031_inst_req_1); -- 
    -- CP-element group 1255 transition  input  bypass 
    -- predecessors 1253 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_4006_to_assign_stmt_4032/type_cast_4031_Sample/ra
      -- 	branch_block_stmt_2042/assign_stmt_4006_to_assign_stmt_4032/type_cast_4031_Sample/$exit
      -- 	branch_block_stmt_2042/assign_stmt_4006_to_assign_stmt_4032/type_cast_4031_sample_completed_
      -- 
    ra_15494_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4031_inst_ack_0, ack => cp_elements(1255)); -- 
    -- CP-element group 1256 fork  transition  place  input  bypass 
    -- predecessors 1254 
    -- successors 2578 2580 
    -- members (11) 
      -- 	branch_block_stmt_2042/assign_stmt_4006_to_assign_stmt_4032__exit__
      -- 	branch_block_stmt_2042/xx_xcritedgex_xi_fdiv32x_xexit
      -- 	branch_block_stmt_2042/assign_stmt_4006_to_assign_stmt_4032/type_cast_4031_Update/$exit
      -- 	branch_block_stmt_2042/assign_stmt_4006_to_assign_stmt_4032/type_cast_4031_Update/ca
      -- 	branch_block_stmt_2042/assign_stmt_4006_to_assign_stmt_4032/$exit
      -- 	branch_block_stmt_2042/assign_stmt_4006_to_assign_stmt_4032/type_cast_4031_update_completed_
      -- 	branch_block_stmt_2042/xx_xcritedgex_xi_fdiv32x_xexit_PhiReq/$entry
      -- 	branch_block_stmt_2042/xx_xcritedgex_xi_fdiv32x_xexit_PhiReq/phi_stmt_4035/$entry
      -- 	branch_block_stmt_2042/xx_xcritedgex_xi_fdiv32x_xexit_PhiReq/phi_stmt_4035/phi_stmt_4035_sources/$entry
      -- 	branch_block_stmt_2042/xx_xcritedgex_xi_fdiv32x_xexit_PhiReq/phi_stmt_4035/phi_stmt_4035_sources/type_cast_4038/$entry
      -- 	branch_block_stmt_2042/xx_xcritedgex_xi_fdiv32x_xexit_PhiReq/phi_stmt_4035/phi_stmt_4035_sources/type_cast_4038/SplitProtocol/$entry
      -- 
    ca_15499_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4031_inst_ack_1, ack => cp_elements(1256)); -- 
    -- CP-element group 1257 fork  transition  bypass 
    -- predecessors 2585 
    -- successors 1258 1259 
    -- members (1) 
      -- 	branch_block_stmt_2042/assign_stmt_4045/$entry
      -- 
    cp_elements(1257) <= cp_elements(2585);
    -- CP-element group 1258 transition  output  bypass 
    -- predecessors 1257 
    -- successors 1260 
    -- members (7) 
      -- 	branch_block_stmt_2042/assign_stmt_4045/WPIPE_out_data_4043_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_4045/R_iNsTr_216_4044_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_4045/R_iNsTr_216_4044_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_4045/WPIPE_out_data_4043_Sample/$entry
      -- 	branch_block_stmt_2042/assign_stmt_4045/R_iNsTr_216_4044_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_4045/R_iNsTr_216_4044_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_4045/WPIPE_out_data_4043_Sample/req
      -- 
    cp_elements(1258) <= cp_elements(1257);
    req_15514_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1258), ack => WPIPE_out_data_4043_inst_req_0); -- 
    -- CP-element group 1259 transition  output  bypass 
    -- predecessors 1257 
    -- successors 1261 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_4045/WPIPE_out_data_4043_Update/$entry
      -- 	branch_block_stmt_2042/assign_stmt_4045/WPIPE_out_data_4043_Update/req
      -- 	branch_block_stmt_2042/assign_stmt_4045/WPIPE_out_data_4043_update_start_
      -- 
    cp_elements(1259) <= cp_elements(1257);
    req_15519_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1259), ack => WPIPE_out_data_4043_inst_req_1); -- 
    -- CP-element group 1260 transition  input  bypass 
    -- predecessors 1258 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_4045/WPIPE_out_data_4043_Sample/ack
      -- 	branch_block_stmt_2042/assign_stmt_4045/WPIPE_out_data_4043_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_4045/WPIPE_out_data_4043_Sample/$exit
      -- 
    ack_15515_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_out_data_4043_inst_ack_0, ack => cp_elements(1260)); -- 
    -- CP-element group 1261 transition  place  input  bypass 
    -- predecessors 1259 
    -- successors 1262 
    -- members (6) 
      -- 	branch_block_stmt_2042/assign_stmt_4045__exit__
      -- 	branch_block_stmt_2042/assign_stmt_4048__entry__
      -- 	branch_block_stmt_2042/assign_stmt_4045/WPIPE_out_data_4043_Update/$exit
      -- 	branch_block_stmt_2042/assign_stmt_4045/WPIPE_out_data_4043_Update/ack
      -- 	branch_block_stmt_2042/assign_stmt_4045/$exit
      -- 	branch_block_stmt_2042/assign_stmt_4045/WPIPE_out_data_4043_update_completed_
      -- 
    ack_15520_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_out_data_4043_inst_ack_1, ack => cp_elements(1261)); -- 
    -- CP-element group 1262 fork  transition  bypass 
    -- predecessors 1261 
    -- successors 1263 1264 
    -- members (1) 
      -- 	branch_block_stmt_2042/assign_stmt_4048/$entry
      -- 
    cp_elements(1262) <= cp_elements(1261);
    -- CP-element group 1263 transition  output  bypass 
    -- predecessors 1262 
    -- successors 1265 
    -- members (7) 
      -- 	branch_block_stmt_2042/assign_stmt_4048/R_iNsTr_81_4047_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_4048/R_iNsTr_81_4047_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_4048/R_iNsTr_81_4047_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_4048/WPIPE_out_data_4046_Sample/req
      -- 	branch_block_stmt_2042/assign_stmt_4048/WPIPE_out_data_4046_Sample/$entry
      -- 	branch_block_stmt_2042/assign_stmt_4048/WPIPE_out_data_4046_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_4048/R_iNsTr_81_4047_update_completed_
      -- 
    cp_elements(1263) <= cp_elements(1262);
    req_15535_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1263), ack => WPIPE_out_data_4046_inst_req_0); -- 
    -- CP-element group 1264 transition  output  bypass 
    -- predecessors 1262 
    -- successors 1266 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_4048/WPIPE_out_data_4046_Update/req
      -- 	branch_block_stmt_2042/assign_stmt_4048/WPIPE_out_data_4046_Update/$entry
      -- 	branch_block_stmt_2042/assign_stmt_4048/WPIPE_out_data_4046_update_start_
      -- 
    cp_elements(1264) <= cp_elements(1262);
    req_15540_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1264), ack => WPIPE_out_data_4046_inst_req_1); -- 
    -- CP-element group 1265 transition  input  bypass 
    -- predecessors 1263 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_4048/WPIPE_out_data_4046_Sample/ack
      -- 	branch_block_stmt_2042/assign_stmt_4048/WPIPE_out_data_4046_Sample/$exit
      -- 	branch_block_stmt_2042/assign_stmt_4048/WPIPE_out_data_4046_sample_completed_
      -- 
    ack_15536_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_out_data_4046_inst_ack_0, ack => cp_elements(1265)); -- 
    -- CP-element group 1266 transition  place  input  bypass 
    -- predecessors 1264 
    -- successors 1267 
    -- members (6) 
      -- 	branch_block_stmt_2042/assign_stmt_4048__exit__
      -- 	branch_block_stmt_2042/assign_stmt_4051__entry__
      -- 	branch_block_stmt_2042/assign_stmt_4048/$exit
      -- 	branch_block_stmt_2042/assign_stmt_4048/WPIPE_out_data_4046_Update/ack
      -- 	branch_block_stmt_2042/assign_stmt_4048/WPIPE_out_data_4046_Update/$exit
      -- 	branch_block_stmt_2042/assign_stmt_4048/WPIPE_out_data_4046_update_completed_
      -- 
    ack_15541_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_out_data_4046_inst_ack_1, ack => cp_elements(1266)); -- 
    -- CP-element group 1267 fork  transition  bypass 
    -- predecessors 1266 
    -- successors 1268 1269 
    -- members (1) 
      -- 	branch_block_stmt_2042/assign_stmt_4051/$entry
      -- 
    cp_elements(1267) <= cp_elements(1266);
    -- CP-element group 1268 transition  output  bypass 
    -- predecessors 1267 
    -- successors 1270 
    -- members (7) 
      -- 	branch_block_stmt_2042/assign_stmt_4051/WPIPE_out_data_4049_Sample/req
      -- 	branch_block_stmt_2042/assign_stmt_4051/WPIPE_out_data_4049_Sample/$entry
      -- 	branch_block_stmt_2042/assign_stmt_4051/WPIPE_out_data_4049_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_4051/R_iNsTr_59_4050_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_4051/R_iNsTr_59_4050_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_4051/R_iNsTr_59_4050_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_4051/R_iNsTr_59_4050_sample_start_
      -- 
    cp_elements(1268) <= cp_elements(1267);
    req_15556_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1268), ack => WPIPE_out_data_4049_inst_req_0); -- 
    -- CP-element group 1269 transition  output  bypass 
    -- predecessors 1267 
    -- successors 1271 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_4051/WPIPE_out_data_4049_Update/req
      -- 	branch_block_stmt_2042/assign_stmt_4051/WPIPE_out_data_4049_Update/$entry
      -- 	branch_block_stmt_2042/assign_stmt_4051/WPIPE_out_data_4049_update_start_
      -- 
    cp_elements(1269) <= cp_elements(1267);
    req_15561_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1269), ack => WPIPE_out_data_4049_inst_req_1); -- 
    -- CP-element group 1270 transition  input  bypass 
    -- predecessors 1268 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_4051/WPIPE_out_data_4049_Sample/ack
      -- 	branch_block_stmt_2042/assign_stmt_4051/WPIPE_out_data_4049_Sample/$exit
      -- 	branch_block_stmt_2042/assign_stmt_4051/WPIPE_out_data_4049_sample_completed_
      -- 
    ack_15557_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_out_data_4049_inst_ack_0, ack => cp_elements(1270)); -- 
    -- CP-element group 1271 transition  place  input  bypass 
    -- predecessors 1269 
    -- successors 1272 
    -- members (6) 
      -- 	branch_block_stmt_2042/assign_stmt_4051__exit__
      -- 	branch_block_stmt_2042/assign_stmt_4054__entry__
      -- 	branch_block_stmt_2042/assign_stmt_4051/WPIPE_out_data_4049_Update/ack
      -- 	branch_block_stmt_2042/assign_stmt_4051/WPIPE_out_data_4049_Update/$exit
      -- 	branch_block_stmt_2042/assign_stmt_4051/WPIPE_out_data_4049_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_4051/$exit
      -- 
    ack_15562_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_out_data_4049_inst_ack_1, ack => cp_elements(1271)); -- 
    -- CP-element group 1272 fork  transition  bypass 
    -- predecessors 1271 
    -- successors 1273 1274 
    -- members (1) 
      -- 	branch_block_stmt_2042/assign_stmt_4054/$entry
      -- 
    cp_elements(1272) <= cp_elements(1271);
    -- CP-element group 1273 transition  output  bypass 
    -- predecessors 1272 
    -- successors 1275 
    -- members (7) 
      -- 	branch_block_stmt_2042/assign_stmt_4054/WPIPE_out_data_4052_Sample/req
      -- 	branch_block_stmt_2042/assign_stmt_4054/WPIPE_out_data_4052_Sample/$entry
      -- 	branch_block_stmt_2042/assign_stmt_4054/WPIPE_out_data_4052_sample_start_
      -- 	branch_block_stmt_2042/assign_stmt_4054/R_iNsTr_42_4053_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_4054/R_iNsTr_42_4053_update_start_
      -- 	branch_block_stmt_2042/assign_stmt_4054/R_iNsTr_42_4053_sample_completed_
      -- 	branch_block_stmt_2042/assign_stmt_4054/R_iNsTr_42_4053_sample_start_
      -- 
    cp_elements(1273) <= cp_elements(1272);
    req_15577_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1273), ack => WPIPE_out_data_4052_inst_req_0); -- 
    -- CP-element group 1274 transition  output  bypass 
    -- predecessors 1272 
    -- successors 1276 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_4054/WPIPE_out_data_4052_Update/req
      -- 	branch_block_stmt_2042/assign_stmt_4054/WPIPE_out_data_4052_Update/$entry
      -- 	branch_block_stmt_2042/assign_stmt_4054/WPIPE_out_data_4052_update_start_
      -- 
    cp_elements(1274) <= cp_elements(1272);
    req_15582_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1274), ack => WPIPE_out_data_4052_inst_req_1); -- 
    -- CP-element group 1275 transition  input  bypass 
    -- predecessors 1273 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_2042/assign_stmt_4054/WPIPE_out_data_4052_Sample/ack
      -- 	branch_block_stmt_2042/assign_stmt_4054/WPIPE_out_data_4052_Sample/$exit
      -- 	branch_block_stmt_2042/assign_stmt_4054/WPIPE_out_data_4052_sample_completed_
      -- 
    ack_15578_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_out_data_4052_inst_ack_0, ack => cp_elements(1275)); -- 
    -- CP-element group 1276 transition  place  input  bypass 
    -- predecessors 1274 
    -- successors 1291 
    -- members (6) 
      -- 	branch_block_stmt_2042/assign_stmt_4054__exit__
      -- 	branch_block_stmt_2042/fdiv32x_xexit_bb_1
      -- 	branch_block_stmt_2042/assign_stmt_4054/WPIPE_out_data_4052_Update/ack
      -- 	branch_block_stmt_2042/assign_stmt_4054/WPIPE_out_data_4052_Update/$exit
      -- 	branch_block_stmt_2042/assign_stmt_4054/WPIPE_out_data_4052_update_completed_
      -- 	branch_block_stmt_2042/assign_stmt_4054/$exit
      -- 
    ack_15583_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_out_data_4052_inst_ack_1, ack => cp_elements(1276)); -- 
    -- CP-element group 1277 fork  transition  bypass 
    -- predecessors 0 
    -- successors 1278 1282 1286 
    -- members (1) 
      -- 	branch_block_stmt_2042/bb_0_bb_1_PhiReq/$entry
      -- 
    cp_elements(1277) <= cp_elements(0);
    -- CP-element group 1278 fork  transition  bypass 
    -- predecessors 1277 
    -- successors 1279 1280 
    -- members (4) 
      -- 	branch_block_stmt_2042/bb_0_bb_1_PhiReq/phi_stmt_2052/$entry
      -- 	branch_block_stmt_2042/bb_0_bb_1_PhiReq/phi_stmt_2052/phi_stmt_2052_sources/$entry
      -- 	branch_block_stmt_2042/bb_0_bb_1_PhiReq/phi_stmt_2052/phi_stmt_2052_sources/type_cast_2058/$entry
      -- 	branch_block_stmt_2042/bb_0_bb_1_PhiReq/phi_stmt_2052/phi_stmt_2052_sources/type_cast_2058/SplitProtocol/$entry
      -- 
    cp_elements(1278) <= cp_elements(1277);
    -- CP-element group 1279 transition  bypass 
    -- predecessors 1278 
    -- successors 1281 
    -- members (4) 
      -- 	branch_block_stmt_2042/bb_0_bb_1_PhiReq/phi_stmt_2052/phi_stmt_2052_sources/type_cast_2058/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_2042/bb_0_bb_1_PhiReq/phi_stmt_2052/phi_stmt_2052_sources/type_cast_2058/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_2042/bb_0_bb_1_PhiReq/phi_stmt_2052/phi_stmt_2052_sources/type_cast_2058/SplitProtocol/Sample/rr
      -- 	branch_block_stmt_2042/bb_0_bb_1_PhiReq/phi_stmt_2052/phi_stmt_2052_sources/type_cast_2058/SplitProtocol/Sample/ra
      -- 
    cp_elements(1279) <= cp_elements(1278);
    -- CP-element group 1280 transition  bypass 
    -- predecessors 1278 
    -- successors 1281 
    -- members (4) 
      -- 	branch_block_stmt_2042/bb_0_bb_1_PhiReq/phi_stmt_2052/phi_stmt_2052_sources/type_cast_2058/SplitProtocol/Update/cr
      -- 	branch_block_stmt_2042/bb_0_bb_1_PhiReq/phi_stmt_2052/phi_stmt_2052_sources/type_cast_2058/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_2042/bb_0_bb_1_PhiReq/phi_stmt_2052/phi_stmt_2052_sources/type_cast_2058/SplitProtocol/Update/ca
      -- 	branch_block_stmt_2042/bb_0_bb_1_PhiReq/phi_stmt_2052/phi_stmt_2052_sources/type_cast_2058/SplitProtocol/Update/$exit
      -- 
    cp_elements(1280) <= cp_elements(1278);
    -- CP-element group 1281 join  transition  output  bypass 
    -- predecessors 1279 1280 
    -- successors 1290 
    -- members (5) 
      -- 	branch_block_stmt_2042/bb_0_bb_1_PhiReq/phi_stmt_2052/$exit
      -- 	branch_block_stmt_2042/bb_0_bb_1_PhiReq/phi_stmt_2052/phi_stmt_2052_req
      -- 	branch_block_stmt_2042/bb_0_bb_1_PhiReq/phi_stmt_2052/phi_stmt_2052_sources/$exit
      -- 	branch_block_stmt_2042/bb_0_bb_1_PhiReq/phi_stmt_2052/phi_stmt_2052_sources/type_cast_2058/$exit
      -- 	branch_block_stmt_2042/bb_0_bb_1_PhiReq/phi_stmt_2052/phi_stmt_2052_sources/type_cast_2058/SplitProtocol/$exit
      -- 
    cp_element_group_1281: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1281"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1279) & cp_elements(1280);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1281), clk => clk, reset => reset); --
    end block;
    phi_stmt_2052_req_15609_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1281), ack => phi_stmt_2052_req_0); -- 
    -- CP-element group 1282 fork  transition  bypass 
    -- predecessors 1277 
    -- successors 1283 1284 
    -- members (4) 
      -- 	branch_block_stmt_2042/bb_0_bb_1_PhiReq/phi_stmt_2045/phi_stmt_2045_sources/type_cast_2051/$entry
      -- 	branch_block_stmt_2042/bb_0_bb_1_PhiReq/phi_stmt_2045/$entry
      -- 	branch_block_stmt_2042/bb_0_bb_1_PhiReq/phi_stmt_2045/phi_stmt_2045_sources/$entry
      -- 	branch_block_stmt_2042/bb_0_bb_1_PhiReq/phi_stmt_2045/phi_stmt_2045_sources/type_cast_2051/SplitProtocol/$entry
      -- 
    cp_elements(1282) <= cp_elements(1277);
    -- CP-element group 1283 transition  bypass 
    -- predecessors 1282 
    -- successors 1285 
    -- members (4) 
      -- 	branch_block_stmt_2042/bb_0_bb_1_PhiReq/phi_stmt_2045/phi_stmt_2045_sources/type_cast_2051/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_2042/bb_0_bb_1_PhiReq/phi_stmt_2045/phi_stmt_2045_sources/type_cast_2051/SplitProtocol/Sample/rr
      -- 	branch_block_stmt_2042/bb_0_bb_1_PhiReq/phi_stmt_2045/phi_stmt_2045_sources/type_cast_2051/SplitProtocol/Sample/ra
      -- 	branch_block_stmt_2042/bb_0_bb_1_PhiReq/phi_stmt_2045/phi_stmt_2045_sources/type_cast_2051/SplitProtocol/Sample/$entry
      -- 
    cp_elements(1283) <= cp_elements(1282);
    -- CP-element group 1284 transition  bypass 
    -- predecessors 1282 
    -- successors 1285 
    -- members (4) 
      -- 	branch_block_stmt_2042/bb_0_bb_1_PhiReq/phi_stmt_2045/phi_stmt_2045_sources/type_cast_2051/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_2042/bb_0_bb_1_PhiReq/phi_stmt_2045/phi_stmt_2045_sources/type_cast_2051/SplitProtocol/Update/ca
      -- 	branch_block_stmt_2042/bb_0_bb_1_PhiReq/phi_stmt_2045/phi_stmt_2045_sources/type_cast_2051/SplitProtocol/Update/cr
      -- 	branch_block_stmt_2042/bb_0_bb_1_PhiReq/phi_stmt_2045/phi_stmt_2045_sources/type_cast_2051/SplitProtocol/Update/$exit
      -- 
    cp_elements(1284) <= cp_elements(1282);
    -- CP-element group 1285 join  transition  output  bypass 
    -- predecessors 1283 1284 
    -- successors 1290 
    -- members (5) 
      -- 	branch_block_stmt_2042/bb_0_bb_1_PhiReq/phi_stmt_2045/phi_stmt_2045_req
      -- 	branch_block_stmt_2042/bb_0_bb_1_PhiReq/phi_stmt_2045/$exit
      -- 	branch_block_stmt_2042/bb_0_bb_1_PhiReq/phi_stmt_2045/phi_stmt_2045_sources/$exit
      -- 	branch_block_stmt_2042/bb_0_bb_1_PhiReq/phi_stmt_2045/phi_stmt_2045_sources/type_cast_2051/SplitProtocol/$exit
      -- 	branch_block_stmt_2042/bb_0_bb_1_PhiReq/phi_stmt_2045/phi_stmt_2045_sources/type_cast_2051/$exit
      -- 
    cp_element_group_1285: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1285"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1283) & cp_elements(1284);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1285), clk => clk, reset => reset); --
    end block;
    phi_stmt_2045_req_15632_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1285), ack => phi_stmt_2045_req_0); -- 
    -- CP-element group 1286 fork  transition  bypass 
    -- predecessors 1277 
    -- successors 1287 1288 
    -- members (4) 
      -- 	branch_block_stmt_2042/bb_0_bb_1_PhiReq/phi_stmt_2059/phi_stmt_2059_sources/type_cast_2065/SplitProtocol/$entry
      -- 	branch_block_stmt_2042/bb_0_bb_1_PhiReq/phi_stmt_2059/phi_stmt_2059_sources/$entry
      -- 	branch_block_stmt_2042/bb_0_bb_1_PhiReq/phi_stmt_2059/$entry
      -- 	branch_block_stmt_2042/bb_0_bb_1_PhiReq/phi_stmt_2059/phi_stmt_2059_sources/type_cast_2065/$entry
      -- 
    cp_elements(1286) <= cp_elements(1277);
    -- CP-element group 1287 transition  bypass 
    -- predecessors 1286 
    -- successors 1289 
    -- members (4) 
      -- 	branch_block_stmt_2042/bb_0_bb_1_PhiReq/phi_stmt_2059/phi_stmt_2059_sources/type_cast_2065/SplitProtocol/Sample/ra
      -- 	branch_block_stmt_2042/bb_0_bb_1_PhiReq/phi_stmt_2059/phi_stmt_2059_sources/type_cast_2065/SplitProtocol/Sample/rr
      -- 	branch_block_stmt_2042/bb_0_bb_1_PhiReq/phi_stmt_2059/phi_stmt_2059_sources/type_cast_2065/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_2042/bb_0_bb_1_PhiReq/phi_stmt_2059/phi_stmt_2059_sources/type_cast_2065/SplitProtocol/Sample/$entry
      -- 
    cp_elements(1287) <= cp_elements(1286);
    -- CP-element group 1288 transition  bypass 
    -- predecessors 1286 
    -- successors 1289 
    -- members (4) 
      -- 	branch_block_stmt_2042/bb_0_bb_1_PhiReq/phi_stmt_2059/phi_stmt_2059_sources/type_cast_2065/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_2042/bb_0_bb_1_PhiReq/phi_stmt_2059/phi_stmt_2059_sources/type_cast_2065/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_2042/bb_0_bb_1_PhiReq/phi_stmt_2059/phi_stmt_2059_sources/type_cast_2065/SplitProtocol/Update/ca
      -- 	branch_block_stmt_2042/bb_0_bb_1_PhiReq/phi_stmt_2059/phi_stmt_2059_sources/type_cast_2065/SplitProtocol/Update/cr
      -- 
    cp_elements(1288) <= cp_elements(1286);
    -- CP-element group 1289 join  transition  output  bypass 
    -- predecessors 1287 1288 
    -- successors 1290 
    -- members (5) 
      -- 	branch_block_stmt_2042/bb_0_bb_1_PhiReq/phi_stmt_2059/$exit
      -- 	branch_block_stmt_2042/bb_0_bb_1_PhiReq/phi_stmt_2059/phi_stmt_2059_sources/type_cast_2065/$exit
      -- 	branch_block_stmt_2042/bb_0_bb_1_PhiReq/phi_stmt_2059/phi_stmt_2059_req
      -- 	branch_block_stmt_2042/bb_0_bb_1_PhiReq/phi_stmt_2059/phi_stmt_2059_sources/$exit
      -- 	branch_block_stmt_2042/bb_0_bb_1_PhiReq/phi_stmt_2059/phi_stmt_2059_sources/type_cast_2065/SplitProtocol/$exit
      -- 
    cp_element_group_1289: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1289"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1287) & cp_elements(1288);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1289), clk => clk, reset => reset); --
    end block;
    phi_stmt_2059_req_15655_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1289), ack => phi_stmt_2059_req_0); -- 
    -- CP-element group 1290 join  transition  bypass 
    -- predecessors 1281 1285 1289 
    -- successors 1311 
    -- members (1) 
      -- 	branch_block_stmt_2042/bb_0_bb_1_PhiReq/$exit
      -- 
    cp_element_group_1290: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1290"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= cp_elements(1281) & cp_elements(1285) & cp_elements(1289);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1290), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1291 fork  transition  bypass 
    -- predecessors 1276 
    -- successors 1292 1298 1304 
    -- members (1) 
      -- 	branch_block_stmt_2042/fdiv32x_xexit_bb_1_PhiReq/$entry
      -- 
    cp_elements(1291) <= cp_elements(1276);
    -- CP-element group 1292 fork  transition  bypass 
    -- predecessors 1291 
    -- successors 1293 1295 
    -- members (4) 
      -- 	branch_block_stmt_2042/fdiv32x_xexit_bb_1_PhiReq/phi_stmt_2052/phi_stmt_2052_sources/type_cast_2058/SplitProtocol/$entry
      -- 	branch_block_stmt_2042/fdiv32x_xexit_bb_1_PhiReq/phi_stmt_2052/$entry
      -- 	branch_block_stmt_2042/fdiv32x_xexit_bb_1_PhiReq/phi_stmt_2052/phi_stmt_2052_sources/type_cast_2058/$entry
      -- 	branch_block_stmt_2042/fdiv32x_xexit_bb_1_PhiReq/phi_stmt_2052/phi_stmt_2052_sources/$entry
      -- 
    cp_elements(1292) <= cp_elements(1291);
    -- CP-element group 1293 transition  output  bypass 
    -- predecessors 1292 
    -- successors 1294 
    -- members (2) 
      -- 	branch_block_stmt_2042/fdiv32x_xexit_bb_1_PhiReq/phi_stmt_2052/phi_stmt_2052_sources/type_cast_2058/SplitProtocol/Sample/rr
      -- 	branch_block_stmt_2042/fdiv32x_xexit_bb_1_PhiReq/phi_stmt_2052/phi_stmt_2052_sources/type_cast_2058/SplitProtocol/Sample/$entry
      -- 
    cp_elements(1293) <= cp_elements(1292);
    rr_15674_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1293), ack => type_cast_2058_inst_req_0); -- 
    -- CP-element group 1294 transition  input  bypass 
    -- predecessors 1293 
    -- successors 1297 
    -- members (2) 
      -- 	branch_block_stmt_2042/fdiv32x_xexit_bb_1_PhiReq/phi_stmt_2052/phi_stmt_2052_sources/type_cast_2058/SplitProtocol/Sample/ra
      -- 	branch_block_stmt_2042/fdiv32x_xexit_bb_1_PhiReq/phi_stmt_2052/phi_stmt_2052_sources/type_cast_2058/SplitProtocol/Sample/$exit
      -- 
    ra_15675_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2058_inst_ack_0, ack => cp_elements(1294)); -- 
    -- CP-element group 1295 transition  output  bypass 
    -- predecessors 1292 
    -- successors 1296 
    -- members (2) 
      -- 	branch_block_stmt_2042/fdiv32x_xexit_bb_1_PhiReq/phi_stmt_2052/phi_stmt_2052_sources/type_cast_2058/SplitProtocol/Update/cr
      -- 	branch_block_stmt_2042/fdiv32x_xexit_bb_1_PhiReq/phi_stmt_2052/phi_stmt_2052_sources/type_cast_2058/SplitProtocol/Update/$entry
      -- 
    cp_elements(1295) <= cp_elements(1292);
    cr_15679_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1295), ack => type_cast_2058_inst_req_1); -- 
    -- CP-element group 1296 transition  input  bypass 
    -- predecessors 1295 
    -- successors 1297 
    -- members (2) 
      -- 	branch_block_stmt_2042/fdiv32x_xexit_bb_1_PhiReq/phi_stmt_2052/phi_stmt_2052_sources/type_cast_2058/SplitProtocol/Update/ca
      -- 	branch_block_stmt_2042/fdiv32x_xexit_bb_1_PhiReq/phi_stmt_2052/phi_stmt_2052_sources/type_cast_2058/SplitProtocol/Update/$exit
      -- 
    ca_15680_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2058_inst_ack_1, ack => cp_elements(1296)); -- 
    -- CP-element group 1297 join  transition  output  bypass 
    -- predecessors 1294 1296 
    -- successors 1310 
    -- members (5) 
      -- 	branch_block_stmt_2042/fdiv32x_xexit_bb_1_PhiReq/phi_stmt_2052/phi_stmt_2052_sources/type_cast_2058/$exit
      -- 	branch_block_stmt_2042/fdiv32x_xexit_bb_1_PhiReq/phi_stmt_2052/phi_stmt_2052_req
      -- 	branch_block_stmt_2042/fdiv32x_xexit_bb_1_PhiReq/phi_stmt_2052/phi_stmt_2052_sources/$exit
      -- 	branch_block_stmt_2042/fdiv32x_xexit_bb_1_PhiReq/phi_stmt_2052/$exit
      -- 	branch_block_stmt_2042/fdiv32x_xexit_bb_1_PhiReq/phi_stmt_2052/phi_stmt_2052_sources/type_cast_2058/SplitProtocol/$exit
      -- 
    cp_element_group_1297: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1297"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1294) & cp_elements(1296);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1297), clk => clk, reset => reset); --
    end block;
    phi_stmt_2052_req_15681_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1297), ack => phi_stmt_2052_req_1); -- 
    -- CP-element group 1298 fork  transition  bypass 
    -- predecessors 1291 
    -- successors 1299 1301 
    -- members (4) 
      -- 	branch_block_stmt_2042/fdiv32x_xexit_bb_1_PhiReq/phi_stmt_2045/phi_stmt_2045_sources/type_cast_2051/SplitProtocol/$entry
      -- 	branch_block_stmt_2042/fdiv32x_xexit_bb_1_PhiReq/phi_stmt_2045/phi_stmt_2045_sources/type_cast_2051/$entry
      -- 	branch_block_stmt_2042/fdiv32x_xexit_bb_1_PhiReq/phi_stmt_2045/phi_stmt_2045_sources/$entry
      -- 	branch_block_stmt_2042/fdiv32x_xexit_bb_1_PhiReq/phi_stmt_2045/$entry
      -- 
    cp_elements(1298) <= cp_elements(1291);
    -- CP-element group 1299 transition  output  bypass 
    -- predecessors 1298 
    -- successors 1300 
    -- members (2) 
      -- 	branch_block_stmt_2042/fdiv32x_xexit_bb_1_PhiReq/phi_stmt_2045/phi_stmt_2045_sources/type_cast_2051/SplitProtocol/Sample/rr
      -- 	branch_block_stmt_2042/fdiv32x_xexit_bb_1_PhiReq/phi_stmt_2045/phi_stmt_2045_sources/type_cast_2051/SplitProtocol/Sample/$entry
      -- 
    cp_elements(1299) <= cp_elements(1298);
    rr_15697_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1299), ack => type_cast_2051_inst_req_0); -- 
    -- CP-element group 1300 transition  input  bypass 
    -- predecessors 1299 
    -- successors 1303 
    -- members (2) 
      -- 	branch_block_stmt_2042/fdiv32x_xexit_bb_1_PhiReq/phi_stmt_2045/phi_stmt_2045_sources/type_cast_2051/SplitProtocol/Sample/ra
      -- 	branch_block_stmt_2042/fdiv32x_xexit_bb_1_PhiReq/phi_stmt_2045/phi_stmt_2045_sources/type_cast_2051/SplitProtocol/Sample/$exit
      -- 
    ra_15698_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2051_inst_ack_0, ack => cp_elements(1300)); -- 
    -- CP-element group 1301 transition  output  bypass 
    -- predecessors 1298 
    -- successors 1302 
    -- members (2) 
      -- 	branch_block_stmt_2042/fdiv32x_xexit_bb_1_PhiReq/phi_stmt_2045/phi_stmt_2045_sources/type_cast_2051/SplitProtocol/Update/cr
      -- 	branch_block_stmt_2042/fdiv32x_xexit_bb_1_PhiReq/phi_stmt_2045/phi_stmt_2045_sources/type_cast_2051/SplitProtocol/Update/$entry
      -- 
    cp_elements(1301) <= cp_elements(1298);
    cr_15702_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1301), ack => type_cast_2051_inst_req_1); -- 
    -- CP-element group 1302 transition  input  bypass 
    -- predecessors 1301 
    -- successors 1303 
    -- members (2) 
      -- 	branch_block_stmt_2042/fdiv32x_xexit_bb_1_PhiReq/phi_stmt_2045/phi_stmt_2045_sources/type_cast_2051/SplitProtocol/Update/ca
      -- 	branch_block_stmt_2042/fdiv32x_xexit_bb_1_PhiReq/phi_stmt_2045/phi_stmt_2045_sources/type_cast_2051/SplitProtocol/Update/$exit
      -- 
    ca_15703_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2051_inst_ack_1, ack => cp_elements(1302)); -- 
    -- CP-element group 1303 join  transition  output  bypass 
    -- predecessors 1300 1302 
    -- successors 1310 
    -- members (5) 
      -- 	branch_block_stmt_2042/fdiv32x_xexit_bb_1_PhiReq/phi_stmt_2045/phi_stmt_2045_req
      -- 	branch_block_stmt_2042/fdiv32x_xexit_bb_1_PhiReq/phi_stmt_2045/phi_stmt_2045_sources/type_cast_2051/SplitProtocol/$exit
      -- 	branch_block_stmt_2042/fdiv32x_xexit_bb_1_PhiReq/phi_stmt_2045/phi_stmt_2045_sources/type_cast_2051/$exit
      -- 	branch_block_stmt_2042/fdiv32x_xexit_bb_1_PhiReq/phi_stmt_2045/phi_stmt_2045_sources/$exit
      -- 	branch_block_stmt_2042/fdiv32x_xexit_bb_1_PhiReq/phi_stmt_2045/$exit
      -- 
    cp_element_group_1303: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1303"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1300) & cp_elements(1302);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1303), clk => clk, reset => reset); --
    end block;
    phi_stmt_2045_req_15704_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1303), ack => phi_stmt_2045_req_1); -- 
    -- CP-element group 1304 fork  transition  bypass 
    -- predecessors 1291 
    -- successors 1305 1307 
    -- members (4) 
      -- 	branch_block_stmt_2042/fdiv32x_xexit_bb_1_PhiReq/phi_stmt_2059/phi_stmt_2059_sources/$entry
      -- 	branch_block_stmt_2042/fdiv32x_xexit_bb_1_PhiReq/phi_stmt_2059/$entry
      -- 	branch_block_stmt_2042/fdiv32x_xexit_bb_1_PhiReq/phi_stmt_2059/phi_stmt_2059_sources/type_cast_2065/SplitProtocol/$entry
      -- 	branch_block_stmt_2042/fdiv32x_xexit_bb_1_PhiReq/phi_stmt_2059/phi_stmt_2059_sources/type_cast_2065/$entry
      -- 
    cp_elements(1304) <= cp_elements(1291);
    -- CP-element group 1305 transition  output  bypass 
    -- predecessors 1304 
    -- successors 1306 
    -- members (2) 
      -- 	branch_block_stmt_2042/fdiv32x_xexit_bb_1_PhiReq/phi_stmt_2059/phi_stmt_2059_sources/type_cast_2065/SplitProtocol/Sample/rr
      -- 	branch_block_stmt_2042/fdiv32x_xexit_bb_1_PhiReq/phi_stmt_2059/phi_stmt_2059_sources/type_cast_2065/SplitProtocol/Sample/$entry
      -- 
    cp_elements(1305) <= cp_elements(1304);
    rr_15720_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1305), ack => type_cast_2065_inst_req_0); -- 
    -- CP-element group 1306 transition  input  bypass 
    -- predecessors 1305 
    -- successors 1309 
    -- members (2) 
      -- 	branch_block_stmt_2042/fdiv32x_xexit_bb_1_PhiReq/phi_stmt_2059/phi_stmt_2059_sources/type_cast_2065/SplitProtocol/Sample/ra
      -- 	branch_block_stmt_2042/fdiv32x_xexit_bb_1_PhiReq/phi_stmt_2059/phi_stmt_2059_sources/type_cast_2065/SplitProtocol/Sample/$exit
      -- 
    ra_15721_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2065_inst_ack_0, ack => cp_elements(1306)); -- 
    -- CP-element group 1307 transition  output  bypass 
    -- predecessors 1304 
    -- successors 1308 
    -- members (2) 
      -- 	branch_block_stmt_2042/fdiv32x_xexit_bb_1_PhiReq/phi_stmt_2059/phi_stmt_2059_sources/type_cast_2065/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_2042/fdiv32x_xexit_bb_1_PhiReq/phi_stmt_2059/phi_stmt_2059_sources/type_cast_2065/SplitProtocol/Update/cr
      -- 
    cp_elements(1307) <= cp_elements(1304);
    cr_15725_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1307), ack => type_cast_2065_inst_req_1); -- 
    -- CP-element group 1308 transition  input  bypass 
    -- predecessors 1307 
    -- successors 1309 
    -- members (2) 
      -- 	branch_block_stmt_2042/fdiv32x_xexit_bb_1_PhiReq/phi_stmt_2059/phi_stmt_2059_sources/type_cast_2065/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_2042/fdiv32x_xexit_bb_1_PhiReq/phi_stmt_2059/phi_stmt_2059_sources/type_cast_2065/SplitProtocol/Update/ca
      -- 
    ca_15726_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2065_inst_ack_1, ack => cp_elements(1308)); -- 
    -- CP-element group 1309 join  transition  output  bypass 
    -- predecessors 1306 1308 
    -- successors 1310 
    -- members (5) 
      -- 	branch_block_stmt_2042/fdiv32x_xexit_bb_1_PhiReq/phi_stmt_2059/phi_stmt_2059_sources/$exit
      -- 	branch_block_stmt_2042/fdiv32x_xexit_bb_1_PhiReq/phi_stmt_2059/$exit
      -- 	branch_block_stmt_2042/fdiv32x_xexit_bb_1_PhiReq/phi_stmt_2059/phi_stmt_2059_req
      -- 	branch_block_stmt_2042/fdiv32x_xexit_bb_1_PhiReq/phi_stmt_2059/phi_stmt_2059_sources/type_cast_2065/SplitProtocol/$exit
      -- 	branch_block_stmt_2042/fdiv32x_xexit_bb_1_PhiReq/phi_stmt_2059/phi_stmt_2059_sources/type_cast_2065/$exit
      -- 
    cp_element_group_1309: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1309"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1306) & cp_elements(1308);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1309), clk => clk, reset => reset); --
    end block;
    phi_stmt_2059_req_15727_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1309), ack => phi_stmt_2059_req_1); -- 
    -- CP-element group 1310 join  transition  bypass 
    -- predecessors 1297 1303 1309 
    -- successors 1311 
    -- members (1) 
      -- 	branch_block_stmt_2042/fdiv32x_xexit_bb_1_PhiReq/$exit
      -- 
    cp_element_group_1310: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1310"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= cp_elements(1297) & cp_elements(1303) & cp_elements(1309);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1310), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1311 merge  place  bypass 
    -- predecessors 1290 1310 
    -- successors 1312 
    -- members (1) 
      -- 	branch_block_stmt_2042/merge_stmt_2044_PhiReqMerge
      -- 
    cp_elements(1311) <= OrReduce(cp_elements(1290) & cp_elements(1310));
    -- CP-element group 1312 fork  transition  bypass 
    -- predecessors 1311 
    -- successors 1313 1314 1315 
    -- members (1) 
      -- 	branch_block_stmt_2042/merge_stmt_2044_PhiAck/$entry
      -- 
    cp_elements(1312) <= cp_elements(1311);
    -- CP-element group 1313 transition  input  bypass 
    -- predecessors 1312 
    -- successors 1316 
    -- members (1) 
      -- 	branch_block_stmt_2042/merge_stmt_2044_PhiAck/phi_stmt_2045_ack
      -- 
    phi_stmt_2045_ack_15732_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2045_ack_0, ack => cp_elements(1313)); -- 
    -- CP-element group 1314 transition  input  bypass 
    -- predecessors 1312 
    -- successors 1316 
    -- members (1) 
      -- 	branch_block_stmt_2042/merge_stmt_2044_PhiAck/phi_stmt_2052_ack
      -- 
    phi_stmt_2052_ack_15733_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2052_ack_0, ack => cp_elements(1314)); -- 
    -- CP-element group 1315 transition  input  bypass 
    -- predecessors 1312 
    -- successors 1316 
    -- members (1) 
      -- 	branch_block_stmt_2042/merge_stmt_2044_PhiAck/phi_stmt_2059_ack
      -- 
    phi_stmt_2059_ack_15734_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2059_ack_0, ack => cp_elements(1315)); -- 
    -- CP-element group 1316 join  transition  bypass 
    -- predecessors 1313 1314 1315 
    -- successors 2 
    -- members (1) 
      -- 	branch_block_stmt_2042/merge_stmt_2044_PhiAck/$exit
      -- 
    cp_element_group_1316: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1316"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= cp_elements(1313) & cp_elements(1314) & cp_elements(1315);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1316), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1317 transition  bypass 
    -- predecessors 127 
    -- successors 1319 
    -- members (4) 
      -- 	branch_block_stmt_2042/bb_1_bb_4_PhiReq/phi_stmt_2134/phi_stmt_2134_sources/type_cast_2137/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_2042/bb_1_bb_4_PhiReq/phi_stmt_2134/phi_stmt_2134_sources/type_cast_2137/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_2042/bb_1_bb_4_PhiReq/phi_stmt_2134/phi_stmt_2134_sources/type_cast_2137/SplitProtocol/Sample/rr
      -- 	branch_block_stmt_2042/bb_1_bb_4_PhiReq/phi_stmt_2134/phi_stmt_2134_sources/type_cast_2137/SplitProtocol/Sample/ra
      -- 
    cp_elements(1317) <= cp_elements(127);
    -- CP-element group 1318 transition  bypass 
    -- predecessors 127 
    -- successors 1319 
    -- members (4) 
      -- 	branch_block_stmt_2042/bb_1_bb_4_PhiReq/phi_stmt_2134/phi_stmt_2134_sources/type_cast_2137/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_2042/bb_1_bb_4_PhiReq/phi_stmt_2134/phi_stmt_2134_sources/type_cast_2137/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_2042/bb_1_bb_4_PhiReq/phi_stmt_2134/phi_stmt_2134_sources/type_cast_2137/SplitProtocol/Update/cr
      -- 	branch_block_stmt_2042/bb_1_bb_4_PhiReq/phi_stmt_2134/phi_stmt_2134_sources/type_cast_2137/SplitProtocol/Update/ca
      -- 
    cp_elements(1318) <= cp_elements(127);
    -- CP-element group 1319 join  transition  output  bypass 
    -- predecessors 1317 1318 
    -- successors 1328 
    -- members (6) 
      -- 	branch_block_stmt_2042/bb_1_bb_4_PhiReq/$exit
      -- 	branch_block_stmt_2042/bb_1_bb_4_PhiReq/phi_stmt_2134/$exit
      -- 	branch_block_stmt_2042/bb_1_bb_4_PhiReq/phi_stmt_2134/phi_stmt_2134_sources/$exit
      -- 	branch_block_stmt_2042/bb_1_bb_4_PhiReq/phi_stmt_2134/phi_stmt_2134_sources/type_cast_2137/$exit
      -- 	branch_block_stmt_2042/bb_1_bb_4_PhiReq/phi_stmt_2134/phi_stmt_2134_sources/type_cast_2137/SplitProtocol/$exit
      -- 	branch_block_stmt_2042/bb_1_bb_4_PhiReq/phi_stmt_2134/phi_stmt_2134_req
      -- 
    cp_element_group_1319: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1319"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1317) & cp_elements(1318);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1319), clk => clk, reset => reset); --
    end block;
    phi_stmt_2134_req_15784_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1319), ack => phi_stmt_2134_req_1); -- 
    -- CP-element group 1320 transition  bypass 
    -- predecessors 139 
    -- successors 1322 
    -- members (4) 
      -- 	branch_block_stmt_2042/bb_2_bb_4_PhiReq/phi_stmt_2134/phi_stmt_2134_sources/type_cast_2137/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_2042/bb_2_bb_4_PhiReq/phi_stmt_2134/phi_stmt_2134_sources/type_cast_2137/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_2042/bb_2_bb_4_PhiReq/phi_stmt_2134/phi_stmt_2134_sources/type_cast_2137/SplitProtocol/Sample/rr
      -- 	branch_block_stmt_2042/bb_2_bb_4_PhiReq/phi_stmt_2134/phi_stmt_2134_sources/type_cast_2137/SplitProtocol/Sample/ra
      -- 
    cp_elements(1320) <= cp_elements(139);
    -- CP-element group 1321 transition  bypass 
    -- predecessors 139 
    -- successors 1322 
    -- members (4) 
      -- 	branch_block_stmt_2042/bb_2_bb_4_PhiReq/phi_stmt_2134/phi_stmt_2134_sources/type_cast_2137/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_2042/bb_2_bb_4_PhiReq/phi_stmt_2134/phi_stmt_2134_sources/type_cast_2137/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_2042/bb_2_bb_4_PhiReq/phi_stmt_2134/phi_stmt_2134_sources/type_cast_2137/SplitProtocol/Update/cr
      -- 	branch_block_stmt_2042/bb_2_bb_4_PhiReq/phi_stmt_2134/phi_stmt_2134_sources/type_cast_2137/SplitProtocol/Update/ca
      -- 
    cp_elements(1321) <= cp_elements(139);
    -- CP-element group 1322 join  transition  output  bypass 
    -- predecessors 1320 1321 
    -- successors 1328 
    -- members (6) 
      -- 	branch_block_stmt_2042/bb_2_bb_4_PhiReq/$exit
      -- 	branch_block_stmt_2042/bb_2_bb_4_PhiReq/phi_stmt_2134/$exit
      -- 	branch_block_stmt_2042/bb_2_bb_4_PhiReq/phi_stmt_2134/phi_stmt_2134_sources/$exit
      -- 	branch_block_stmt_2042/bb_2_bb_4_PhiReq/phi_stmt_2134/phi_stmt_2134_sources/type_cast_2137/$exit
      -- 	branch_block_stmt_2042/bb_2_bb_4_PhiReq/phi_stmt_2134/phi_stmt_2134_sources/type_cast_2137/SplitProtocol/$exit
      -- 	branch_block_stmt_2042/bb_2_bb_4_PhiReq/phi_stmt_2134/phi_stmt_2134_req
      -- 
    cp_element_group_1322: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1322"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1320) & cp_elements(1321);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1322), clk => clk, reset => reset); --
    end block;
    phi_stmt_2134_req_15810_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1322), ack => phi_stmt_2134_req_2); -- 
    -- CP-element group 1323 transition  output  bypass 
    -- predecessors 4 
    -- successors 1324 
    -- members (2) 
      -- 	branch_block_stmt_2042/bb_3_bb_4_PhiReq/phi_stmt_2134/phi_stmt_2134_sources/type_cast_2137/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_2042/bb_3_bb_4_PhiReq/phi_stmt_2134/phi_stmt_2134_sources/type_cast_2137/SplitProtocol/Sample/rr
      -- 
    cp_elements(1323) <= cp_elements(4);
    rr_15829_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1323), ack => type_cast_2137_inst_req_0); -- 
    -- CP-element group 1324 transition  input  bypass 
    -- predecessors 1323 
    -- successors 1327 
    -- members (2) 
      -- 	branch_block_stmt_2042/bb_3_bb_4_PhiReq/phi_stmt_2134/phi_stmt_2134_sources/type_cast_2137/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_2042/bb_3_bb_4_PhiReq/phi_stmt_2134/phi_stmt_2134_sources/type_cast_2137/SplitProtocol/Sample/ra
      -- 
    ra_15830_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2137_inst_ack_0, ack => cp_elements(1324)); -- 
    -- CP-element group 1325 transition  output  bypass 
    -- predecessors 4 
    -- successors 1326 
    -- members (2) 
      -- 	branch_block_stmt_2042/bb_3_bb_4_PhiReq/phi_stmt_2134/phi_stmt_2134_sources/type_cast_2137/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_2042/bb_3_bb_4_PhiReq/phi_stmt_2134/phi_stmt_2134_sources/type_cast_2137/SplitProtocol/Update/cr
      -- 
    cp_elements(1325) <= cp_elements(4);
    cr_15834_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1325), ack => type_cast_2137_inst_req_1); -- 
    -- CP-element group 1326 transition  input  bypass 
    -- predecessors 1325 
    -- successors 1327 
    -- members (2) 
      -- 	branch_block_stmt_2042/bb_3_bb_4_PhiReq/phi_stmt_2134/phi_stmt_2134_sources/type_cast_2137/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_2042/bb_3_bb_4_PhiReq/phi_stmt_2134/phi_stmt_2134_sources/type_cast_2137/SplitProtocol/Update/ca
      -- 
    ca_15835_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2137_inst_ack_1, ack => cp_elements(1326)); -- 
    -- CP-element group 1327 join  transition  output  bypass 
    -- predecessors 1324 1326 
    -- successors 1328 
    -- members (6) 
      -- 	branch_block_stmt_2042/bb_3_bb_4_PhiReq/$exit
      -- 	branch_block_stmt_2042/bb_3_bb_4_PhiReq/phi_stmt_2134/$exit
      -- 	branch_block_stmt_2042/bb_3_bb_4_PhiReq/phi_stmt_2134/phi_stmt_2134_sources/$exit
      -- 	branch_block_stmt_2042/bb_3_bb_4_PhiReq/phi_stmt_2134/phi_stmt_2134_sources/type_cast_2137/$exit
      -- 	branch_block_stmt_2042/bb_3_bb_4_PhiReq/phi_stmt_2134/phi_stmt_2134_sources/type_cast_2137/SplitProtocol/$exit
      -- 	branch_block_stmt_2042/bb_3_bb_4_PhiReq/phi_stmt_2134/phi_stmt_2134_req
      -- 
    cp_element_group_1327: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1327"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1324) & cp_elements(1326);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1327), clk => clk, reset => reset); --
    end block;
    phi_stmt_2134_req_15836_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1327), ack => phi_stmt_2134_req_0); -- 
    -- CP-element group 1328 merge  place  bypass 
    -- predecessors 1319 1322 1327 
    -- successors 1329 
    -- members (1) 
      -- 	branch_block_stmt_2042/merge_stmt_2133_PhiReqMerge
      -- 
    cp_elements(1328) <= OrReduce(cp_elements(1319) & cp_elements(1322) & cp_elements(1327));
    -- CP-element group 1329 transition  bypass 
    -- predecessors 1328 
    -- successors 1330 
    -- members (1) 
      -- 	branch_block_stmt_2042/merge_stmt_2133_PhiAck/$entry
      -- 
    cp_elements(1329) <= cp_elements(1328);
    -- CP-element group 1330 transition  place  input  bypass 
    -- predecessors 1329 
    -- successors 142 
    -- members (4) 
      -- 	branch_block_stmt_2042/merge_stmt_2133__exit__
      -- 	branch_block_stmt_2042/assign_stmt_2150_to_assign_stmt_2161__entry__
      -- 	branch_block_stmt_2042/merge_stmt_2133_PhiAck/$exit
      -- 	branch_block_stmt_2042/merge_stmt_2133_PhiAck/phi_stmt_2134_ack
      -- 
    phi_stmt_2134_ack_15841_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2134_ack_0, ack => cp_elements(1330)); -- 
    -- CP-element group 1331 transition  bypass 
    -- predecessors 159 
    -- successors 1333 
    -- members (4) 
      -- 	branch_block_stmt_2042/bb_4_bb_7_PhiReq/phi_stmt_2190/phi_stmt_2190_sources/type_cast_2193/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_2042/bb_4_bb_7_PhiReq/phi_stmt_2190/phi_stmt_2190_sources/type_cast_2193/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_2042/bb_4_bb_7_PhiReq/phi_stmt_2190/phi_stmt_2190_sources/type_cast_2193/SplitProtocol/Sample/rr
      -- 	branch_block_stmt_2042/bb_4_bb_7_PhiReq/phi_stmt_2190/phi_stmt_2190_sources/type_cast_2193/SplitProtocol/Sample/ra
      -- 
    cp_elements(1331) <= cp_elements(159);
    -- CP-element group 1332 transition  bypass 
    -- predecessors 159 
    -- successors 1333 
    -- members (4) 
      -- 	branch_block_stmt_2042/bb_4_bb_7_PhiReq/phi_stmt_2190/phi_stmt_2190_sources/type_cast_2193/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_2042/bb_4_bb_7_PhiReq/phi_stmt_2190/phi_stmt_2190_sources/type_cast_2193/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_2042/bb_4_bb_7_PhiReq/phi_stmt_2190/phi_stmt_2190_sources/type_cast_2193/SplitProtocol/Update/cr
      -- 	branch_block_stmt_2042/bb_4_bb_7_PhiReq/phi_stmt_2190/phi_stmt_2190_sources/type_cast_2193/SplitProtocol/Update/ca
      -- 
    cp_elements(1332) <= cp_elements(159);
    -- CP-element group 1333 join  transition  output  bypass 
    -- predecessors 1331 1332 
    -- successors 1342 
    -- members (6) 
      -- 	branch_block_stmt_2042/bb_4_bb_7_PhiReq/$exit
      -- 	branch_block_stmt_2042/bb_4_bb_7_PhiReq/phi_stmt_2190/$exit
      -- 	branch_block_stmt_2042/bb_4_bb_7_PhiReq/phi_stmt_2190/phi_stmt_2190_sources/$exit
      -- 	branch_block_stmt_2042/bb_4_bb_7_PhiReq/phi_stmt_2190/phi_stmt_2190_sources/type_cast_2193/$exit
      -- 	branch_block_stmt_2042/bb_4_bb_7_PhiReq/phi_stmt_2190/phi_stmt_2190_sources/type_cast_2193/SplitProtocol/$exit
      -- 	branch_block_stmt_2042/bb_4_bb_7_PhiReq/phi_stmt_2190/phi_stmt_2190_req
      -- 
    cp_element_group_1333: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1333"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1331) & cp_elements(1332);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1333), clk => clk, reset => reset); --
    end block;
    phi_stmt_2190_req_15891_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1333), ack => phi_stmt_2190_req_1); -- 
    -- CP-element group 1334 transition  bypass 
    -- predecessors 171 
    -- successors 1336 
    -- members (4) 
      -- 	branch_block_stmt_2042/bb_5_bb_7_PhiReq/phi_stmt_2190/phi_stmt_2190_sources/type_cast_2193/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_2042/bb_5_bb_7_PhiReq/phi_stmt_2190/phi_stmt_2190_sources/type_cast_2193/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_2042/bb_5_bb_7_PhiReq/phi_stmt_2190/phi_stmt_2190_sources/type_cast_2193/SplitProtocol/Sample/rr
      -- 	branch_block_stmt_2042/bb_5_bb_7_PhiReq/phi_stmt_2190/phi_stmt_2190_sources/type_cast_2193/SplitProtocol/Sample/ra
      -- 
    cp_elements(1334) <= cp_elements(171);
    -- CP-element group 1335 transition  bypass 
    -- predecessors 171 
    -- successors 1336 
    -- members (4) 
      -- 	branch_block_stmt_2042/bb_5_bb_7_PhiReq/phi_stmt_2190/phi_stmt_2190_sources/type_cast_2193/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_2042/bb_5_bb_7_PhiReq/phi_stmt_2190/phi_stmt_2190_sources/type_cast_2193/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_2042/bb_5_bb_7_PhiReq/phi_stmt_2190/phi_stmt_2190_sources/type_cast_2193/SplitProtocol/Update/cr
      -- 	branch_block_stmt_2042/bb_5_bb_7_PhiReq/phi_stmt_2190/phi_stmt_2190_sources/type_cast_2193/SplitProtocol/Update/ca
      -- 
    cp_elements(1335) <= cp_elements(171);
    -- CP-element group 1336 join  transition  output  bypass 
    -- predecessors 1334 1335 
    -- successors 1342 
    -- members (6) 
      -- 	branch_block_stmt_2042/bb_5_bb_7_PhiReq/$exit
      -- 	branch_block_stmt_2042/bb_5_bb_7_PhiReq/phi_stmt_2190/$exit
      -- 	branch_block_stmt_2042/bb_5_bb_7_PhiReq/phi_stmt_2190/phi_stmt_2190_sources/$exit
      -- 	branch_block_stmt_2042/bb_5_bb_7_PhiReq/phi_stmt_2190/phi_stmt_2190_sources/type_cast_2193/$exit
      -- 	branch_block_stmt_2042/bb_5_bb_7_PhiReq/phi_stmt_2190/phi_stmt_2190_sources/type_cast_2193/SplitProtocol/$exit
      -- 	branch_block_stmt_2042/bb_5_bb_7_PhiReq/phi_stmt_2190/phi_stmt_2190_req
      -- 
    cp_element_group_1336: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1336"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1334) & cp_elements(1335);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1336), clk => clk, reset => reset); --
    end block;
    phi_stmt_2190_req_15917_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1336), ack => phi_stmt_2190_req_2); -- 
    -- CP-element group 1337 transition  output  bypass 
    -- predecessors 178 
    -- successors 1338 
    -- members (2) 
      -- 	branch_block_stmt_2042/bb_6_bb_7_PhiReq/phi_stmt_2190/phi_stmt_2190_sources/type_cast_2193/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_2042/bb_6_bb_7_PhiReq/phi_stmt_2190/phi_stmt_2190_sources/type_cast_2193/SplitProtocol/Sample/rr
      -- 
    cp_elements(1337) <= cp_elements(178);
    rr_15936_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1337), ack => type_cast_2193_inst_req_0); -- 
    -- CP-element group 1338 transition  input  bypass 
    -- predecessors 1337 
    -- successors 1341 
    -- members (2) 
      -- 	branch_block_stmt_2042/bb_6_bb_7_PhiReq/phi_stmt_2190/phi_stmt_2190_sources/type_cast_2193/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_2042/bb_6_bb_7_PhiReq/phi_stmt_2190/phi_stmt_2190_sources/type_cast_2193/SplitProtocol/Sample/ra
      -- 
    ra_15937_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2193_inst_ack_0, ack => cp_elements(1338)); -- 
    -- CP-element group 1339 transition  output  bypass 
    -- predecessors 178 
    -- successors 1340 
    -- members (2) 
      -- 	branch_block_stmt_2042/bb_6_bb_7_PhiReq/phi_stmt_2190/phi_stmt_2190_sources/type_cast_2193/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_2042/bb_6_bb_7_PhiReq/phi_stmt_2190/phi_stmt_2190_sources/type_cast_2193/SplitProtocol/Update/cr
      -- 
    cp_elements(1339) <= cp_elements(178);
    cr_15941_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1339), ack => type_cast_2193_inst_req_1); -- 
    -- CP-element group 1340 transition  input  bypass 
    -- predecessors 1339 
    -- successors 1341 
    -- members (2) 
      -- 	branch_block_stmt_2042/bb_6_bb_7_PhiReq/phi_stmt_2190/phi_stmt_2190_sources/type_cast_2193/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_2042/bb_6_bb_7_PhiReq/phi_stmt_2190/phi_stmt_2190_sources/type_cast_2193/SplitProtocol/Update/ca
      -- 
    ca_15942_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2193_inst_ack_1, ack => cp_elements(1340)); -- 
    -- CP-element group 1341 join  transition  output  bypass 
    -- predecessors 1338 1340 
    -- successors 1342 
    -- members (6) 
      -- 	branch_block_stmt_2042/bb_6_bb_7_PhiReq/$exit
      -- 	branch_block_stmt_2042/bb_6_bb_7_PhiReq/phi_stmt_2190/$exit
      -- 	branch_block_stmt_2042/bb_6_bb_7_PhiReq/phi_stmt_2190/phi_stmt_2190_sources/$exit
      -- 	branch_block_stmt_2042/bb_6_bb_7_PhiReq/phi_stmt_2190/phi_stmt_2190_sources/type_cast_2193/$exit
      -- 	branch_block_stmt_2042/bb_6_bb_7_PhiReq/phi_stmt_2190/phi_stmt_2190_sources/type_cast_2193/SplitProtocol/$exit
      -- 	branch_block_stmt_2042/bb_6_bb_7_PhiReq/phi_stmt_2190/phi_stmt_2190_req
      -- 
    cp_element_group_1341: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1341"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1338) & cp_elements(1340);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1341), clk => clk, reset => reset); --
    end block;
    phi_stmt_2190_req_15943_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1341), ack => phi_stmt_2190_req_0); -- 
    -- CP-element group 1342 merge  place  bypass 
    -- predecessors 1333 1336 1341 
    -- successors 1343 
    -- members (1) 
      -- 	branch_block_stmt_2042/merge_stmt_2189_PhiReqMerge
      -- 
    cp_elements(1342) <= OrReduce(cp_elements(1333) & cp_elements(1336) & cp_elements(1341));
    -- CP-element group 1343 transition  bypass 
    -- predecessors 1342 
    -- successors 1344 
    -- members (1) 
      -- 	branch_block_stmt_2042/merge_stmt_2189_PhiAck/$entry
      -- 
    cp_elements(1343) <= cp_elements(1342);
    -- CP-element group 1344 transition  place  input  bypass 
    -- predecessors 1343 
    -- successors 179 
    -- members (4) 
      -- 	branch_block_stmt_2042/merge_stmt_2189__exit__
      -- 	branch_block_stmt_2042/assign_stmt_2204_to_assign_stmt_2210__entry__
      -- 	branch_block_stmt_2042/merge_stmt_2189_PhiAck/$exit
      -- 	branch_block_stmt_2042/merge_stmt_2189_PhiAck/phi_stmt_2190_ack
      -- 
    phi_stmt_2190_ack_15948_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2190_ack_0, ack => cp_elements(1344)); -- 
    -- CP-element group 1345 fork  transition  bypass 
    -- predecessors 239 
    -- successors 1346 1347 
    -- members (2) 
      -- 	branch_block_stmt_2042/bb_11_bb_13_PhiReq/phi_stmt_2304/phi_stmt_2304_sources/type_cast_2307/$entry
      -- 	branch_block_stmt_2042/bb_11_bb_13_PhiReq/phi_stmt_2304/phi_stmt_2304_sources/type_cast_2307/SplitProtocol/$entry
      -- 
    cp_elements(1345) <= cp_elements(239);
    -- CP-element group 1346 transition  bypass 
    -- predecessors 1345 
    -- successors 1348 
    -- members (4) 
      -- 	branch_block_stmt_2042/bb_11_bb_13_PhiReq/phi_stmt_2304/phi_stmt_2304_sources/type_cast_2307/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_2042/bb_11_bb_13_PhiReq/phi_stmt_2304/phi_stmt_2304_sources/type_cast_2307/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_2042/bb_11_bb_13_PhiReq/phi_stmt_2304/phi_stmt_2304_sources/type_cast_2307/SplitProtocol/Sample/rr
      -- 	branch_block_stmt_2042/bb_11_bb_13_PhiReq/phi_stmt_2304/phi_stmt_2304_sources/type_cast_2307/SplitProtocol/Sample/ra
      -- 
    cp_elements(1346) <= cp_elements(1345);
    -- CP-element group 1347 transition  bypass 
    -- predecessors 1345 
    -- successors 1348 
    -- members (4) 
      -- 	branch_block_stmt_2042/bb_11_bb_13_PhiReq/phi_stmt_2304/phi_stmt_2304_sources/type_cast_2307/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_2042/bb_11_bb_13_PhiReq/phi_stmt_2304/phi_stmt_2304_sources/type_cast_2307/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_2042/bb_11_bb_13_PhiReq/phi_stmt_2304/phi_stmt_2304_sources/type_cast_2307/SplitProtocol/Update/cr
      -- 	branch_block_stmt_2042/bb_11_bb_13_PhiReq/phi_stmt_2304/phi_stmt_2304_sources/type_cast_2307/SplitProtocol/Update/ca
      -- 
    cp_elements(1347) <= cp_elements(1345);
    -- CP-element group 1348 join  transition  bypass 
    -- predecessors 1346 1347 
    -- successors 1359 
    -- members (2) 
      -- 	branch_block_stmt_2042/bb_11_bb_13_PhiReq/phi_stmt_2304/phi_stmt_2304_sources/type_cast_2307/$exit
      -- 	branch_block_stmt_2042/bb_11_bb_13_PhiReq/phi_stmt_2304/phi_stmt_2304_sources/type_cast_2307/SplitProtocol/$exit
      -- 
    cp_element_group_1348: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1348"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1346) & cp_elements(1347);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1348), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1349 fork  transition  bypass 
    -- predecessors 239 
    -- successors 1350 1352 
    -- members (2) 
      -- 	branch_block_stmt_2042/bb_11_bb_13_PhiReq/phi_stmt_2304/phi_stmt_2304_sources/type_cast_2309/$entry
      -- 	branch_block_stmt_2042/bb_11_bb_13_PhiReq/phi_stmt_2304/phi_stmt_2304_sources/type_cast_2309/SplitProtocol/$entry
      -- 
    cp_elements(1349) <= cp_elements(239);
    -- CP-element group 1350 transition  output  bypass 
    -- predecessors 1349 
    -- successors 1351 
    -- members (2) 
      -- 	branch_block_stmt_2042/bb_11_bb_13_PhiReq/phi_stmt_2304/phi_stmt_2304_sources/type_cast_2309/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_2042/bb_11_bb_13_PhiReq/phi_stmt_2304/phi_stmt_2304_sources/type_cast_2309/SplitProtocol/Sample/rr
      -- 
    cp_elements(1350) <= cp_elements(1349);
    rr_16035_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1350), ack => type_cast_2309_inst_req_0); -- 
    -- CP-element group 1351 transition  input  bypass 
    -- predecessors 1350 
    -- successors 1354 
    -- members (2) 
      -- 	branch_block_stmt_2042/bb_11_bb_13_PhiReq/phi_stmt_2304/phi_stmt_2304_sources/type_cast_2309/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_2042/bb_11_bb_13_PhiReq/phi_stmt_2304/phi_stmt_2304_sources/type_cast_2309/SplitProtocol/Sample/ra
      -- 
    ra_16036_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2309_inst_ack_0, ack => cp_elements(1351)); -- 
    -- CP-element group 1352 transition  output  bypass 
    -- predecessors 1349 
    -- successors 1353 
    -- members (2) 
      -- 	branch_block_stmt_2042/bb_11_bb_13_PhiReq/phi_stmt_2304/phi_stmt_2304_sources/type_cast_2309/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_2042/bb_11_bb_13_PhiReq/phi_stmt_2304/phi_stmt_2304_sources/type_cast_2309/SplitProtocol/Update/cr
      -- 
    cp_elements(1352) <= cp_elements(1349);
    cr_16040_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1352), ack => type_cast_2309_inst_req_1); -- 
    -- CP-element group 1353 transition  input  bypass 
    -- predecessors 1352 
    -- successors 1354 
    -- members (2) 
      -- 	branch_block_stmt_2042/bb_11_bb_13_PhiReq/phi_stmt_2304/phi_stmt_2304_sources/type_cast_2309/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_2042/bb_11_bb_13_PhiReq/phi_stmt_2304/phi_stmt_2304_sources/type_cast_2309/SplitProtocol/Update/ca
      -- 
    ca_16041_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2309_inst_ack_1, ack => cp_elements(1353)); -- 
    -- CP-element group 1354 join  transition  bypass 
    -- predecessors 1351 1353 
    -- successors 1359 
    -- members (2) 
      -- 	branch_block_stmt_2042/bb_11_bb_13_PhiReq/phi_stmt_2304/phi_stmt_2304_sources/type_cast_2309/$exit
      -- 	branch_block_stmt_2042/bb_11_bb_13_PhiReq/phi_stmt_2304/phi_stmt_2304_sources/type_cast_2309/SplitProtocol/$exit
      -- 
    cp_element_group_1354: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1354"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1351) & cp_elements(1353);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1354), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1355 fork  transition  bypass 
    -- predecessors 239 
    -- successors 1356 1357 
    -- members (2) 
      -- 	branch_block_stmt_2042/bb_11_bb_13_PhiReq/phi_stmt_2304/phi_stmt_2304_sources/type_cast_2311/$entry
      -- 	branch_block_stmt_2042/bb_11_bb_13_PhiReq/phi_stmt_2304/phi_stmt_2304_sources/type_cast_2311/SplitProtocol/$entry
      -- 
    cp_elements(1355) <= cp_elements(239);
    -- CP-element group 1356 transition  bypass 
    -- predecessors 1355 
    -- successors 1358 
    -- members (4) 
      -- 	branch_block_stmt_2042/bb_11_bb_13_PhiReq/phi_stmt_2304/phi_stmt_2304_sources/type_cast_2311/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_2042/bb_11_bb_13_PhiReq/phi_stmt_2304/phi_stmt_2304_sources/type_cast_2311/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_2042/bb_11_bb_13_PhiReq/phi_stmt_2304/phi_stmt_2304_sources/type_cast_2311/SplitProtocol/Sample/rr
      -- 	branch_block_stmt_2042/bb_11_bb_13_PhiReq/phi_stmt_2304/phi_stmt_2304_sources/type_cast_2311/SplitProtocol/Sample/ra
      -- 
    cp_elements(1356) <= cp_elements(1355);
    -- CP-element group 1357 transition  bypass 
    -- predecessors 1355 
    -- successors 1358 
    -- members (4) 
      -- 	branch_block_stmt_2042/bb_11_bb_13_PhiReq/phi_stmt_2304/phi_stmt_2304_sources/type_cast_2311/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_2042/bb_11_bb_13_PhiReq/phi_stmt_2304/phi_stmt_2304_sources/type_cast_2311/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_2042/bb_11_bb_13_PhiReq/phi_stmt_2304/phi_stmt_2304_sources/type_cast_2311/SplitProtocol/Update/cr
      -- 	branch_block_stmt_2042/bb_11_bb_13_PhiReq/phi_stmt_2304/phi_stmt_2304_sources/type_cast_2311/SplitProtocol/Update/ca
      -- 
    cp_elements(1357) <= cp_elements(1355);
    -- CP-element group 1358 join  transition  bypass 
    -- predecessors 1356 1357 
    -- successors 1359 
    -- members (2) 
      -- 	branch_block_stmt_2042/bb_11_bb_13_PhiReq/phi_stmt_2304/phi_stmt_2304_sources/type_cast_2311/$exit
      -- 	branch_block_stmt_2042/bb_11_bb_13_PhiReq/phi_stmt_2304/phi_stmt_2304_sources/type_cast_2311/SplitProtocol/$exit
      -- 
    cp_element_group_1358: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1358"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1356) & cp_elements(1357);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1358), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1359 join  transition  output  bypass 
    -- predecessors 1348 1354 1358 
    -- successors 1403 
    -- members (4) 
      -- 	branch_block_stmt_2042/bb_11_bb_13_PhiReq/$exit
      -- 	branch_block_stmt_2042/bb_11_bb_13_PhiReq/phi_stmt_2304/$exit
      -- 	branch_block_stmt_2042/bb_11_bb_13_PhiReq/phi_stmt_2304/phi_stmt_2304_sources/$exit
      -- 	branch_block_stmt_2042/bb_11_bb_13_PhiReq/phi_stmt_2304/phi_stmt_2304_req
      -- 
    cp_element_group_1359: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1359"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= cp_elements(1348) & cp_elements(1354) & cp_elements(1358);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1359), clk => clk, reset => reset); --
    end block;
    phi_stmt_2304_req_16058_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1359), ack => phi_stmt_2304_req_1); -- 
    -- CP-element group 1360 fork  transition  bypass 
    -- predecessors 250 
    -- successors 1361 1362 
    -- members (2) 
      -- 	branch_block_stmt_2042/bb_12_bb_13_PhiReq/phi_stmt_2304/phi_stmt_2304_sources/type_cast_2307/$entry
      -- 	branch_block_stmt_2042/bb_12_bb_13_PhiReq/phi_stmt_2304/phi_stmt_2304_sources/type_cast_2307/SplitProtocol/$entry
      -- 
    cp_elements(1360) <= cp_elements(250);
    -- CP-element group 1361 transition  bypass 
    -- predecessors 1360 
    -- successors 1363 
    -- members (4) 
      -- 	branch_block_stmt_2042/bb_12_bb_13_PhiReq/phi_stmt_2304/phi_stmt_2304_sources/type_cast_2307/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_2042/bb_12_bb_13_PhiReq/phi_stmt_2304/phi_stmt_2304_sources/type_cast_2307/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_2042/bb_12_bb_13_PhiReq/phi_stmt_2304/phi_stmt_2304_sources/type_cast_2307/SplitProtocol/Sample/rr
      -- 	branch_block_stmt_2042/bb_12_bb_13_PhiReq/phi_stmt_2304/phi_stmt_2304_sources/type_cast_2307/SplitProtocol/Sample/ra
      -- 
    cp_elements(1361) <= cp_elements(1360);
    -- CP-element group 1362 transition  bypass 
    -- predecessors 1360 
    -- successors 1363 
    -- members (4) 
      -- 	branch_block_stmt_2042/bb_12_bb_13_PhiReq/phi_stmt_2304/phi_stmt_2304_sources/type_cast_2307/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_2042/bb_12_bb_13_PhiReq/phi_stmt_2304/phi_stmt_2304_sources/type_cast_2307/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_2042/bb_12_bb_13_PhiReq/phi_stmt_2304/phi_stmt_2304_sources/type_cast_2307/SplitProtocol/Update/cr
      -- 	branch_block_stmt_2042/bb_12_bb_13_PhiReq/phi_stmt_2304/phi_stmt_2304_sources/type_cast_2307/SplitProtocol/Update/ca
      -- 
    cp_elements(1362) <= cp_elements(1360);
    -- CP-element group 1363 join  transition  bypass 
    -- predecessors 1361 1362 
    -- successors 1374 
    -- members (2) 
      -- 	branch_block_stmt_2042/bb_12_bb_13_PhiReq/phi_stmt_2304/phi_stmt_2304_sources/type_cast_2307/$exit
      -- 	branch_block_stmt_2042/bb_12_bb_13_PhiReq/phi_stmt_2304/phi_stmt_2304_sources/type_cast_2307/SplitProtocol/$exit
      -- 
    cp_element_group_1363: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1363"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1361) & cp_elements(1362);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1363), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1364 fork  transition  bypass 
    -- predecessors 250 
    -- successors 1365 1366 
    -- members (2) 
      -- 	branch_block_stmt_2042/bb_12_bb_13_PhiReq/phi_stmt_2304/phi_stmt_2304_sources/type_cast_2309/$entry
      -- 	branch_block_stmt_2042/bb_12_bb_13_PhiReq/phi_stmt_2304/phi_stmt_2304_sources/type_cast_2309/SplitProtocol/$entry
      -- 
    cp_elements(1364) <= cp_elements(250);
    -- CP-element group 1365 transition  bypass 
    -- predecessors 1364 
    -- successors 1367 
    -- members (4) 
      -- 	branch_block_stmt_2042/bb_12_bb_13_PhiReq/phi_stmt_2304/phi_stmt_2304_sources/type_cast_2309/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_2042/bb_12_bb_13_PhiReq/phi_stmt_2304/phi_stmt_2304_sources/type_cast_2309/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_2042/bb_12_bb_13_PhiReq/phi_stmt_2304/phi_stmt_2304_sources/type_cast_2309/SplitProtocol/Sample/rr
      -- 	branch_block_stmt_2042/bb_12_bb_13_PhiReq/phi_stmt_2304/phi_stmt_2304_sources/type_cast_2309/SplitProtocol/Sample/ra
      -- 
    cp_elements(1365) <= cp_elements(1364);
    -- CP-element group 1366 transition  bypass 
    -- predecessors 1364 
    -- successors 1367 
    -- members (4) 
      -- 	branch_block_stmt_2042/bb_12_bb_13_PhiReq/phi_stmt_2304/phi_stmt_2304_sources/type_cast_2309/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_2042/bb_12_bb_13_PhiReq/phi_stmt_2304/phi_stmt_2304_sources/type_cast_2309/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_2042/bb_12_bb_13_PhiReq/phi_stmt_2304/phi_stmt_2304_sources/type_cast_2309/SplitProtocol/Update/cr
      -- 	branch_block_stmt_2042/bb_12_bb_13_PhiReq/phi_stmt_2304/phi_stmt_2304_sources/type_cast_2309/SplitProtocol/Update/ca
      -- 
    cp_elements(1366) <= cp_elements(1364);
    -- CP-element group 1367 join  transition  bypass 
    -- predecessors 1365 1366 
    -- successors 1374 
    -- members (2) 
      -- 	branch_block_stmt_2042/bb_12_bb_13_PhiReq/phi_stmt_2304/phi_stmt_2304_sources/type_cast_2309/$exit
      -- 	branch_block_stmt_2042/bb_12_bb_13_PhiReq/phi_stmt_2304/phi_stmt_2304_sources/type_cast_2309/SplitProtocol/$exit
      -- 
    cp_element_group_1367: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1367"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1365) & cp_elements(1366);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1367), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1368 fork  transition  bypass 
    -- predecessors 250 
    -- successors 1369 1371 
    -- members (2) 
      -- 	branch_block_stmt_2042/bb_12_bb_13_PhiReq/phi_stmt_2304/phi_stmt_2304_sources/type_cast_2311/$entry
      -- 	branch_block_stmt_2042/bb_12_bb_13_PhiReq/phi_stmt_2304/phi_stmt_2304_sources/type_cast_2311/SplitProtocol/$entry
      -- 
    cp_elements(1368) <= cp_elements(250);
    -- CP-element group 1369 transition  output  bypass 
    -- predecessors 1368 
    -- successors 1370 
    -- members (2) 
      -- 	branch_block_stmt_2042/bb_12_bb_13_PhiReq/phi_stmt_2304/phi_stmt_2304_sources/type_cast_2311/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_2042/bb_12_bb_13_PhiReq/phi_stmt_2304/phi_stmt_2304_sources/type_cast_2311/SplitProtocol/Sample/rr
      -- 
    cp_elements(1369) <= cp_elements(1368);
    rr_16109_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1369), ack => type_cast_2311_inst_req_0); -- 
    -- CP-element group 1370 transition  input  bypass 
    -- predecessors 1369 
    -- successors 1373 
    -- members (2) 
      -- 	branch_block_stmt_2042/bb_12_bb_13_PhiReq/phi_stmt_2304/phi_stmt_2304_sources/type_cast_2311/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_2042/bb_12_bb_13_PhiReq/phi_stmt_2304/phi_stmt_2304_sources/type_cast_2311/SplitProtocol/Sample/ra
      -- 
    ra_16110_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2311_inst_ack_0, ack => cp_elements(1370)); -- 
    -- CP-element group 1371 transition  output  bypass 
    -- predecessors 1368 
    -- successors 1372 
    -- members (2) 
      -- 	branch_block_stmt_2042/bb_12_bb_13_PhiReq/phi_stmt_2304/phi_stmt_2304_sources/type_cast_2311/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_2042/bb_12_bb_13_PhiReq/phi_stmt_2304/phi_stmt_2304_sources/type_cast_2311/SplitProtocol/Update/cr
      -- 
    cp_elements(1371) <= cp_elements(1368);
    cr_16114_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1371), ack => type_cast_2311_inst_req_1); -- 
    -- CP-element group 1372 transition  input  bypass 
    -- predecessors 1371 
    -- successors 1373 
    -- members (2) 
      -- 	branch_block_stmt_2042/bb_12_bb_13_PhiReq/phi_stmt_2304/phi_stmt_2304_sources/type_cast_2311/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_2042/bb_12_bb_13_PhiReq/phi_stmt_2304/phi_stmt_2304_sources/type_cast_2311/SplitProtocol/Update/ca
      -- 
    ca_16115_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2311_inst_ack_1, ack => cp_elements(1372)); -- 
    -- CP-element group 1373 join  transition  bypass 
    -- predecessors 1370 1372 
    -- successors 1374 
    -- members (2) 
      -- 	branch_block_stmt_2042/bb_12_bb_13_PhiReq/phi_stmt_2304/phi_stmt_2304_sources/type_cast_2311/$exit
      -- 	branch_block_stmt_2042/bb_12_bb_13_PhiReq/phi_stmt_2304/phi_stmt_2304_sources/type_cast_2311/SplitProtocol/$exit
      -- 
    cp_element_group_1373: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1373"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1370) & cp_elements(1372);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1373), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1374 join  transition  output  bypass 
    -- predecessors 1363 1367 1373 
    -- successors 1403 
    -- members (4) 
      -- 	branch_block_stmt_2042/bb_12_bb_13_PhiReq/$exit
      -- 	branch_block_stmt_2042/bb_12_bb_13_PhiReq/phi_stmt_2304/$exit
      -- 	branch_block_stmt_2042/bb_12_bb_13_PhiReq/phi_stmt_2304/phi_stmt_2304_sources/$exit
      -- 	branch_block_stmt_2042/bb_12_bb_13_PhiReq/phi_stmt_2304/phi_stmt_2304_req
      -- 
    cp_element_group_1374: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1374"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= cp_elements(1363) & cp_elements(1367) & cp_elements(1373);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1374), clk => clk, reset => reset); --
    end block;
    phi_stmt_2304_req_16116_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1374), ack => phi_stmt_2304_req_2); -- 
    -- CP-element group 1375 fork  transition  bypass 
    -- predecessors 193 
    -- successors 1376 1377 
    -- members (2) 
      -- 	branch_block_stmt_2042/bb_7_bb_13_PhiReq/phi_stmt_2304/phi_stmt_2304_sources/type_cast_2307/$entry
      -- 	branch_block_stmt_2042/bb_7_bb_13_PhiReq/phi_stmt_2304/phi_stmt_2304_sources/type_cast_2307/SplitProtocol/$entry
      -- 
    cp_elements(1375) <= cp_elements(193);
    -- CP-element group 1376 transition  bypass 
    -- predecessors 1375 
    -- successors 1378 
    -- members (4) 
      -- 	branch_block_stmt_2042/bb_7_bb_13_PhiReq/phi_stmt_2304/phi_stmt_2304_sources/type_cast_2307/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_2042/bb_7_bb_13_PhiReq/phi_stmt_2304/phi_stmt_2304_sources/type_cast_2307/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_2042/bb_7_bb_13_PhiReq/phi_stmt_2304/phi_stmt_2304_sources/type_cast_2307/SplitProtocol/Sample/rr
      -- 	branch_block_stmt_2042/bb_7_bb_13_PhiReq/phi_stmt_2304/phi_stmt_2304_sources/type_cast_2307/SplitProtocol/Sample/ra
      -- 
    cp_elements(1376) <= cp_elements(1375);
    -- CP-element group 1377 transition  bypass 
    -- predecessors 1375 
    -- successors 1378 
    -- members (4) 
      -- 	branch_block_stmt_2042/bb_7_bb_13_PhiReq/phi_stmt_2304/phi_stmt_2304_sources/type_cast_2307/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_2042/bb_7_bb_13_PhiReq/phi_stmt_2304/phi_stmt_2304_sources/type_cast_2307/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_2042/bb_7_bb_13_PhiReq/phi_stmt_2304/phi_stmt_2304_sources/type_cast_2307/SplitProtocol/Update/cr
      -- 	branch_block_stmt_2042/bb_7_bb_13_PhiReq/phi_stmt_2304/phi_stmt_2304_sources/type_cast_2307/SplitProtocol/Update/ca
      -- 
    cp_elements(1377) <= cp_elements(1375);
    -- CP-element group 1378 join  transition  bypass 
    -- predecessors 1376 1377 
    -- successors 1387 
    -- members (2) 
      -- 	branch_block_stmt_2042/bb_7_bb_13_PhiReq/phi_stmt_2304/phi_stmt_2304_sources/type_cast_2307/$exit
      -- 	branch_block_stmt_2042/bb_7_bb_13_PhiReq/phi_stmt_2304/phi_stmt_2304_sources/type_cast_2307/SplitProtocol/$exit
      -- 
    cp_element_group_1378: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1378"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1376) & cp_elements(1377);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1378), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1379 fork  transition  bypass 
    -- predecessors 193 
    -- successors 1380 1381 
    -- members (2) 
      -- 	branch_block_stmt_2042/bb_7_bb_13_PhiReq/phi_stmt_2304/phi_stmt_2304_sources/type_cast_2309/$entry
      -- 	branch_block_stmt_2042/bb_7_bb_13_PhiReq/phi_stmt_2304/phi_stmt_2304_sources/type_cast_2309/SplitProtocol/$entry
      -- 
    cp_elements(1379) <= cp_elements(193);
    -- CP-element group 1380 transition  bypass 
    -- predecessors 1379 
    -- successors 1382 
    -- members (4) 
      -- 	branch_block_stmt_2042/bb_7_bb_13_PhiReq/phi_stmt_2304/phi_stmt_2304_sources/type_cast_2309/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_2042/bb_7_bb_13_PhiReq/phi_stmt_2304/phi_stmt_2304_sources/type_cast_2309/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_2042/bb_7_bb_13_PhiReq/phi_stmt_2304/phi_stmt_2304_sources/type_cast_2309/SplitProtocol/Sample/rr
      -- 	branch_block_stmt_2042/bb_7_bb_13_PhiReq/phi_stmt_2304/phi_stmt_2304_sources/type_cast_2309/SplitProtocol/Sample/ra
      -- 
    cp_elements(1380) <= cp_elements(1379);
    -- CP-element group 1381 transition  bypass 
    -- predecessors 1379 
    -- successors 1382 
    -- members (4) 
      -- 	branch_block_stmt_2042/bb_7_bb_13_PhiReq/phi_stmt_2304/phi_stmt_2304_sources/type_cast_2309/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_2042/bb_7_bb_13_PhiReq/phi_stmt_2304/phi_stmt_2304_sources/type_cast_2309/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_2042/bb_7_bb_13_PhiReq/phi_stmt_2304/phi_stmt_2304_sources/type_cast_2309/SplitProtocol/Update/cr
      -- 	branch_block_stmt_2042/bb_7_bb_13_PhiReq/phi_stmt_2304/phi_stmt_2304_sources/type_cast_2309/SplitProtocol/Update/ca
      -- 
    cp_elements(1381) <= cp_elements(1379);
    -- CP-element group 1382 join  transition  bypass 
    -- predecessors 1380 1381 
    -- successors 1387 
    -- members (2) 
      -- 	branch_block_stmt_2042/bb_7_bb_13_PhiReq/phi_stmt_2304/phi_stmt_2304_sources/type_cast_2309/$exit
      -- 	branch_block_stmt_2042/bb_7_bb_13_PhiReq/phi_stmt_2304/phi_stmt_2304_sources/type_cast_2309/SplitProtocol/$exit
      -- 
    cp_element_group_1382: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1382"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1380) & cp_elements(1381);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1382), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1383 fork  transition  bypass 
    -- predecessors 193 
    -- successors 1384 1385 
    -- members (2) 
      -- 	branch_block_stmt_2042/bb_7_bb_13_PhiReq/phi_stmt_2304/phi_stmt_2304_sources/type_cast_2311/$entry
      -- 	branch_block_stmt_2042/bb_7_bb_13_PhiReq/phi_stmt_2304/phi_stmt_2304_sources/type_cast_2311/SplitProtocol/$entry
      -- 
    cp_elements(1383) <= cp_elements(193);
    -- CP-element group 1384 transition  bypass 
    -- predecessors 1383 
    -- successors 1386 
    -- members (4) 
      -- 	branch_block_stmt_2042/bb_7_bb_13_PhiReq/phi_stmt_2304/phi_stmt_2304_sources/type_cast_2311/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_2042/bb_7_bb_13_PhiReq/phi_stmt_2304/phi_stmt_2304_sources/type_cast_2311/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_2042/bb_7_bb_13_PhiReq/phi_stmt_2304/phi_stmt_2304_sources/type_cast_2311/SplitProtocol/Sample/rr
      -- 	branch_block_stmt_2042/bb_7_bb_13_PhiReq/phi_stmt_2304/phi_stmt_2304_sources/type_cast_2311/SplitProtocol/Sample/ra
      -- 
    cp_elements(1384) <= cp_elements(1383);
    -- CP-element group 1385 transition  bypass 
    -- predecessors 1383 
    -- successors 1386 
    -- members (4) 
      -- 	branch_block_stmt_2042/bb_7_bb_13_PhiReq/phi_stmt_2304/phi_stmt_2304_sources/type_cast_2311/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_2042/bb_7_bb_13_PhiReq/phi_stmt_2304/phi_stmt_2304_sources/type_cast_2311/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_2042/bb_7_bb_13_PhiReq/phi_stmt_2304/phi_stmt_2304_sources/type_cast_2311/SplitProtocol/Update/cr
      -- 	branch_block_stmt_2042/bb_7_bb_13_PhiReq/phi_stmt_2304/phi_stmt_2304_sources/type_cast_2311/SplitProtocol/Update/ca
      -- 
    cp_elements(1385) <= cp_elements(1383);
    -- CP-element group 1386 join  transition  bypass 
    -- predecessors 1384 1385 
    -- successors 1387 
    -- members (2) 
      -- 	branch_block_stmt_2042/bb_7_bb_13_PhiReq/phi_stmt_2304/phi_stmt_2304_sources/type_cast_2311/$exit
      -- 	branch_block_stmt_2042/bb_7_bb_13_PhiReq/phi_stmt_2304/phi_stmt_2304_sources/type_cast_2311/SplitProtocol/$exit
      -- 
    cp_element_group_1386: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1386"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1384) & cp_elements(1385);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1386), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1387 join  transition  output  bypass 
    -- predecessors 1378 1382 1386 
    -- successors 1403 
    -- members (4) 
      -- 	branch_block_stmt_2042/bb_7_bb_13_PhiReq/$exit
      -- 	branch_block_stmt_2042/bb_7_bb_13_PhiReq/phi_stmt_2304/$exit
      -- 	branch_block_stmt_2042/bb_7_bb_13_PhiReq/phi_stmt_2304/phi_stmt_2304_sources/$exit
      -- 	branch_block_stmt_2042/bb_7_bb_13_PhiReq/phi_stmt_2304/phi_stmt_2304_req
      -- 
    cp_element_group_1387: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1387"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= cp_elements(1378) & cp_elements(1382) & cp_elements(1386);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1387), clk => clk, reset => reset); --
    end block;
    phi_stmt_2304_req_16174_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1387), ack => phi_stmt_2304_req_3); -- 
    -- CP-element group 1388 fork  transition  bypass 
    -- predecessors 216 
    -- successors 1389 1391 
    -- members (2) 
      -- 	branch_block_stmt_2042/bb_9_bb_13_PhiReq/phi_stmt_2304/phi_stmt_2304_sources/type_cast_2307/$entry
      -- 	branch_block_stmt_2042/bb_9_bb_13_PhiReq/phi_stmt_2304/phi_stmt_2304_sources/type_cast_2307/SplitProtocol/$entry
      -- 
    cp_elements(1388) <= cp_elements(216);
    -- CP-element group 1389 transition  output  bypass 
    -- predecessors 1388 
    -- successors 1390 
    -- members (2) 
      -- 	branch_block_stmt_2042/bb_9_bb_13_PhiReq/phi_stmt_2304/phi_stmt_2304_sources/type_cast_2307/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_2042/bb_9_bb_13_PhiReq/phi_stmt_2304/phi_stmt_2304_sources/type_cast_2307/SplitProtocol/Sample/rr
      -- 
    cp_elements(1389) <= cp_elements(1388);
    rr_16193_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1389), ack => type_cast_2307_inst_req_0); -- 
    -- CP-element group 1390 transition  input  bypass 
    -- predecessors 1389 
    -- successors 1393 
    -- members (2) 
      -- 	branch_block_stmt_2042/bb_9_bb_13_PhiReq/phi_stmt_2304/phi_stmt_2304_sources/type_cast_2307/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_2042/bb_9_bb_13_PhiReq/phi_stmt_2304/phi_stmt_2304_sources/type_cast_2307/SplitProtocol/Sample/ra
      -- 
    ra_16194_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2307_inst_ack_0, ack => cp_elements(1390)); -- 
    -- CP-element group 1391 transition  output  bypass 
    -- predecessors 1388 
    -- successors 1392 
    -- members (2) 
      -- 	branch_block_stmt_2042/bb_9_bb_13_PhiReq/phi_stmt_2304/phi_stmt_2304_sources/type_cast_2307/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_2042/bb_9_bb_13_PhiReq/phi_stmt_2304/phi_stmt_2304_sources/type_cast_2307/SplitProtocol/Update/cr
      -- 
    cp_elements(1391) <= cp_elements(1388);
    cr_16198_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1391), ack => type_cast_2307_inst_req_1); -- 
    -- CP-element group 1392 transition  input  bypass 
    -- predecessors 1391 
    -- successors 1393 
    -- members (2) 
      -- 	branch_block_stmt_2042/bb_9_bb_13_PhiReq/phi_stmt_2304/phi_stmt_2304_sources/type_cast_2307/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_2042/bb_9_bb_13_PhiReq/phi_stmt_2304/phi_stmt_2304_sources/type_cast_2307/SplitProtocol/Update/ca
      -- 
    ca_16199_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2307_inst_ack_1, ack => cp_elements(1392)); -- 
    -- CP-element group 1393 join  transition  bypass 
    -- predecessors 1390 1392 
    -- successors 1402 
    -- members (2) 
      -- 	branch_block_stmt_2042/bb_9_bb_13_PhiReq/phi_stmt_2304/phi_stmt_2304_sources/type_cast_2307/$exit
      -- 	branch_block_stmt_2042/bb_9_bb_13_PhiReq/phi_stmt_2304/phi_stmt_2304_sources/type_cast_2307/SplitProtocol/$exit
      -- 
    cp_element_group_1393: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1393"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1390) & cp_elements(1392);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1393), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1394 fork  transition  bypass 
    -- predecessors 216 
    -- successors 1395 1396 
    -- members (2) 
      -- 	branch_block_stmt_2042/bb_9_bb_13_PhiReq/phi_stmt_2304/phi_stmt_2304_sources/type_cast_2309/$entry
      -- 	branch_block_stmt_2042/bb_9_bb_13_PhiReq/phi_stmt_2304/phi_stmt_2304_sources/type_cast_2309/SplitProtocol/$entry
      -- 
    cp_elements(1394) <= cp_elements(216);
    -- CP-element group 1395 transition  bypass 
    -- predecessors 1394 
    -- successors 1397 
    -- members (4) 
      -- 	branch_block_stmt_2042/bb_9_bb_13_PhiReq/phi_stmt_2304/phi_stmt_2304_sources/type_cast_2309/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_2042/bb_9_bb_13_PhiReq/phi_stmt_2304/phi_stmt_2304_sources/type_cast_2309/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_2042/bb_9_bb_13_PhiReq/phi_stmt_2304/phi_stmt_2304_sources/type_cast_2309/SplitProtocol/Sample/rr
      -- 	branch_block_stmt_2042/bb_9_bb_13_PhiReq/phi_stmt_2304/phi_stmt_2304_sources/type_cast_2309/SplitProtocol/Sample/ra
      -- 
    cp_elements(1395) <= cp_elements(1394);
    -- CP-element group 1396 transition  bypass 
    -- predecessors 1394 
    -- successors 1397 
    -- members (4) 
      -- 	branch_block_stmt_2042/bb_9_bb_13_PhiReq/phi_stmt_2304/phi_stmt_2304_sources/type_cast_2309/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_2042/bb_9_bb_13_PhiReq/phi_stmt_2304/phi_stmt_2304_sources/type_cast_2309/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_2042/bb_9_bb_13_PhiReq/phi_stmt_2304/phi_stmt_2304_sources/type_cast_2309/SplitProtocol/Update/cr
      -- 	branch_block_stmt_2042/bb_9_bb_13_PhiReq/phi_stmt_2304/phi_stmt_2304_sources/type_cast_2309/SplitProtocol/Update/ca
      -- 
    cp_elements(1396) <= cp_elements(1394);
    -- CP-element group 1397 join  transition  bypass 
    -- predecessors 1395 1396 
    -- successors 1402 
    -- members (2) 
      -- 	branch_block_stmt_2042/bb_9_bb_13_PhiReq/phi_stmt_2304/phi_stmt_2304_sources/type_cast_2309/$exit
      -- 	branch_block_stmt_2042/bb_9_bb_13_PhiReq/phi_stmt_2304/phi_stmt_2304_sources/type_cast_2309/SplitProtocol/$exit
      -- 
    cp_element_group_1397: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1397"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1395) & cp_elements(1396);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1397), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1398 fork  transition  bypass 
    -- predecessors 216 
    -- successors 1399 1400 
    -- members (2) 
      -- 	branch_block_stmt_2042/bb_9_bb_13_PhiReq/phi_stmt_2304/phi_stmt_2304_sources/type_cast_2311/$entry
      -- 	branch_block_stmt_2042/bb_9_bb_13_PhiReq/phi_stmt_2304/phi_stmt_2304_sources/type_cast_2311/SplitProtocol/$entry
      -- 
    cp_elements(1398) <= cp_elements(216);
    -- CP-element group 1399 transition  bypass 
    -- predecessors 1398 
    -- successors 1401 
    -- members (4) 
      -- 	branch_block_stmt_2042/bb_9_bb_13_PhiReq/phi_stmt_2304/phi_stmt_2304_sources/type_cast_2311/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_2042/bb_9_bb_13_PhiReq/phi_stmt_2304/phi_stmt_2304_sources/type_cast_2311/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_2042/bb_9_bb_13_PhiReq/phi_stmt_2304/phi_stmt_2304_sources/type_cast_2311/SplitProtocol/Sample/rr
      -- 	branch_block_stmt_2042/bb_9_bb_13_PhiReq/phi_stmt_2304/phi_stmt_2304_sources/type_cast_2311/SplitProtocol/Sample/ra
      -- 
    cp_elements(1399) <= cp_elements(1398);
    -- CP-element group 1400 transition  bypass 
    -- predecessors 1398 
    -- successors 1401 
    -- members (4) 
      -- 	branch_block_stmt_2042/bb_9_bb_13_PhiReq/phi_stmt_2304/phi_stmt_2304_sources/type_cast_2311/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_2042/bb_9_bb_13_PhiReq/phi_stmt_2304/phi_stmt_2304_sources/type_cast_2311/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_2042/bb_9_bb_13_PhiReq/phi_stmt_2304/phi_stmt_2304_sources/type_cast_2311/SplitProtocol/Update/cr
      -- 	branch_block_stmt_2042/bb_9_bb_13_PhiReq/phi_stmt_2304/phi_stmt_2304_sources/type_cast_2311/SplitProtocol/Update/ca
      -- 
    cp_elements(1400) <= cp_elements(1398);
    -- CP-element group 1401 join  transition  bypass 
    -- predecessors 1399 1400 
    -- successors 1402 
    -- members (2) 
      -- 	branch_block_stmt_2042/bb_9_bb_13_PhiReq/phi_stmt_2304/phi_stmt_2304_sources/type_cast_2311/$exit
      -- 	branch_block_stmt_2042/bb_9_bb_13_PhiReq/phi_stmt_2304/phi_stmt_2304_sources/type_cast_2311/SplitProtocol/$exit
      -- 
    cp_element_group_1401: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1401"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1399) & cp_elements(1400);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1401), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1402 join  transition  output  bypass 
    -- predecessors 1393 1397 1401 
    -- successors 1403 
    -- members (4) 
      -- 	branch_block_stmt_2042/bb_9_bb_13_PhiReq/$exit
      -- 	branch_block_stmt_2042/bb_9_bb_13_PhiReq/phi_stmt_2304/$exit
      -- 	branch_block_stmt_2042/bb_9_bb_13_PhiReq/phi_stmt_2304/phi_stmt_2304_sources/$exit
      -- 	branch_block_stmt_2042/bb_9_bb_13_PhiReq/phi_stmt_2304/phi_stmt_2304_req
      -- 
    cp_element_group_1402: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1402"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= cp_elements(1393) & cp_elements(1397) & cp_elements(1401);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1402), clk => clk, reset => reset); --
    end block;
    phi_stmt_2304_req_16232_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1402), ack => phi_stmt_2304_req_0); -- 
    -- CP-element group 1403 merge  place  bypass 
    -- predecessors 1359 1374 1387 1402 
    -- successors 1404 
    -- members (1) 
      -- 	branch_block_stmt_2042/merge_stmt_2303_PhiReqMerge
      -- 
    cp_elements(1403) <= OrReduce(cp_elements(1359) & cp_elements(1374) & cp_elements(1387) & cp_elements(1402));
    -- CP-element group 1404 transition  bypass 
    -- predecessors 1403 
    -- successors 1405 
    -- members (1) 
      -- 	branch_block_stmt_2042/merge_stmt_2303_PhiAck/$entry
      -- 
    cp_elements(1404) <= cp_elements(1403);
    -- CP-element group 1405 transition  place  input  bypass 
    -- predecessors 1404 
    -- successors 251 
    -- members (4) 
      -- 	branch_block_stmt_2042/merge_stmt_2303__exit__
      -- 	branch_block_stmt_2042/assign_stmt_2321_to_assign_stmt_2342__entry__
      -- 	branch_block_stmt_2042/merge_stmt_2303_PhiAck/$exit
      -- 	branch_block_stmt_2042/merge_stmt_2303_PhiAck/phi_stmt_2304_ack
      -- 
    phi_stmt_2304_ack_16237_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2304_ack_0, ack => cp_elements(1405)); -- 
    -- CP-element group 1406 fork  transition  bypass 
    -- predecessors 290 
    -- successors 1407 1419 
    -- members (1) 
      -- 	branch_block_stmt_2042/bb_14_bbx_xnph7x_xix_xix_xi33_PhiReq/$entry
      -- 
    cp_elements(1406) <= cp_elements(290);
    -- CP-element group 1407 fork  transition  bypass 
    -- predecessors 1406 
    -- successors 1408 1412 
    -- members (2) 
      -- 	branch_block_stmt_2042/bb_14_bbx_xnph7x_xix_xix_xi33_PhiReq/phi_stmt_2370/$entry
      -- 	branch_block_stmt_2042/bb_14_bbx_xnph7x_xix_xix_xi33_PhiReq/phi_stmt_2370/phi_stmt_2370_sources/$entry
      -- 
    cp_elements(1407) <= cp_elements(1406);
    -- CP-element group 1408 fork  transition  bypass 
    -- predecessors 1407 
    -- successors 1409 1410 
    -- members (2) 
      -- 	branch_block_stmt_2042/bb_14_bbx_xnph7x_xix_xix_xi33_PhiReq/phi_stmt_2370/phi_stmt_2370_sources/type_cast_2373/$entry
      -- 	branch_block_stmt_2042/bb_14_bbx_xnph7x_xix_xix_xi33_PhiReq/phi_stmt_2370/phi_stmt_2370_sources/type_cast_2373/SplitProtocol/$entry
      -- 
    cp_elements(1408) <= cp_elements(1407);
    -- CP-element group 1409 transition  bypass 
    -- predecessors 1408 
    -- successors 1411 
    -- members (4) 
      -- 	branch_block_stmt_2042/bb_14_bbx_xnph7x_xix_xix_xi33_PhiReq/phi_stmt_2370/phi_stmt_2370_sources/type_cast_2373/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_2042/bb_14_bbx_xnph7x_xix_xix_xi33_PhiReq/phi_stmt_2370/phi_stmt_2370_sources/type_cast_2373/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_2042/bb_14_bbx_xnph7x_xix_xix_xi33_PhiReq/phi_stmt_2370/phi_stmt_2370_sources/type_cast_2373/SplitProtocol/Sample/rr
      -- 	branch_block_stmt_2042/bb_14_bbx_xnph7x_xix_xix_xi33_PhiReq/phi_stmt_2370/phi_stmt_2370_sources/type_cast_2373/SplitProtocol/Sample/ra
      -- 
    cp_elements(1409) <= cp_elements(1408);
    -- CP-element group 1410 transition  bypass 
    -- predecessors 1408 
    -- successors 1411 
    -- members (4) 
      -- 	branch_block_stmt_2042/bb_14_bbx_xnph7x_xix_xix_xi33_PhiReq/phi_stmt_2370/phi_stmt_2370_sources/type_cast_2373/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_2042/bb_14_bbx_xnph7x_xix_xix_xi33_PhiReq/phi_stmt_2370/phi_stmt_2370_sources/type_cast_2373/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_2042/bb_14_bbx_xnph7x_xix_xix_xi33_PhiReq/phi_stmt_2370/phi_stmt_2370_sources/type_cast_2373/SplitProtocol/Update/cr
      -- 	branch_block_stmt_2042/bb_14_bbx_xnph7x_xix_xix_xi33_PhiReq/phi_stmt_2370/phi_stmt_2370_sources/type_cast_2373/SplitProtocol/Update/ca
      -- 
    cp_elements(1410) <= cp_elements(1408);
    -- CP-element group 1411 join  transition  bypass 
    -- predecessors 1409 1410 
    -- successors 1418 
    -- members (2) 
      -- 	branch_block_stmt_2042/bb_14_bbx_xnph7x_xix_xix_xi33_PhiReq/phi_stmt_2370/phi_stmt_2370_sources/type_cast_2373/$exit
      -- 	branch_block_stmt_2042/bb_14_bbx_xnph7x_xix_xix_xi33_PhiReq/phi_stmt_2370/phi_stmt_2370_sources/type_cast_2373/SplitProtocol/$exit
      -- 
    cp_element_group_1411: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1411"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1409) & cp_elements(1410);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1411), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1412 fork  transition  bypass 
    -- predecessors 1407 
    -- successors 1413 1415 
    -- members (2) 
      -- 	branch_block_stmt_2042/bb_14_bbx_xnph7x_xix_xix_xi33_PhiReq/phi_stmt_2370/phi_stmt_2370_sources/type_cast_2375/$entry
      -- 	branch_block_stmt_2042/bb_14_bbx_xnph7x_xix_xix_xi33_PhiReq/phi_stmt_2370/phi_stmt_2370_sources/type_cast_2375/SplitProtocol/$entry
      -- 
    cp_elements(1412) <= cp_elements(1407);
    -- CP-element group 1413 transition  output  bypass 
    -- predecessors 1412 
    -- successors 1414 
    -- members (2) 
      -- 	branch_block_stmt_2042/bb_14_bbx_xnph7x_xix_xix_xi33_PhiReq/phi_stmt_2370/phi_stmt_2370_sources/type_cast_2375/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_2042/bb_14_bbx_xnph7x_xix_xix_xi33_PhiReq/phi_stmt_2370/phi_stmt_2370_sources/type_cast_2375/SplitProtocol/Sample/rr
      -- 
    cp_elements(1413) <= cp_elements(1412);
    rr_16284_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1413), ack => type_cast_2375_inst_req_0); -- 
    -- CP-element group 1414 transition  input  bypass 
    -- predecessors 1413 
    -- successors 1417 
    -- members (2) 
      -- 	branch_block_stmt_2042/bb_14_bbx_xnph7x_xix_xix_xi33_PhiReq/phi_stmt_2370/phi_stmt_2370_sources/type_cast_2375/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_2042/bb_14_bbx_xnph7x_xix_xix_xi33_PhiReq/phi_stmt_2370/phi_stmt_2370_sources/type_cast_2375/SplitProtocol/Sample/ra
      -- 
    ra_16285_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2375_inst_ack_0, ack => cp_elements(1414)); -- 
    -- CP-element group 1415 transition  output  bypass 
    -- predecessors 1412 
    -- successors 1416 
    -- members (2) 
      -- 	branch_block_stmt_2042/bb_14_bbx_xnph7x_xix_xix_xi33_PhiReq/phi_stmt_2370/phi_stmt_2370_sources/type_cast_2375/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_2042/bb_14_bbx_xnph7x_xix_xix_xi33_PhiReq/phi_stmt_2370/phi_stmt_2370_sources/type_cast_2375/SplitProtocol/Update/cr
      -- 
    cp_elements(1415) <= cp_elements(1412);
    cr_16289_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1415), ack => type_cast_2375_inst_req_1); -- 
    -- CP-element group 1416 transition  input  bypass 
    -- predecessors 1415 
    -- successors 1417 
    -- members (2) 
      -- 	branch_block_stmt_2042/bb_14_bbx_xnph7x_xix_xix_xi33_PhiReq/phi_stmt_2370/phi_stmt_2370_sources/type_cast_2375/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_2042/bb_14_bbx_xnph7x_xix_xix_xi33_PhiReq/phi_stmt_2370/phi_stmt_2370_sources/type_cast_2375/SplitProtocol/Update/ca
      -- 
    ca_16290_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2375_inst_ack_1, ack => cp_elements(1416)); -- 
    -- CP-element group 1417 join  transition  bypass 
    -- predecessors 1414 1416 
    -- successors 1418 
    -- members (2) 
      -- 	branch_block_stmt_2042/bb_14_bbx_xnph7x_xix_xix_xi33_PhiReq/phi_stmt_2370/phi_stmt_2370_sources/type_cast_2375/$exit
      -- 	branch_block_stmt_2042/bb_14_bbx_xnph7x_xix_xix_xi33_PhiReq/phi_stmt_2370/phi_stmt_2370_sources/type_cast_2375/SplitProtocol/$exit
      -- 
    cp_element_group_1417: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1417"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1414) & cp_elements(1416);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1417), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1418 join  transition  output  bypass 
    -- predecessors 1411 1417 
    -- successors 1423 
    -- members (3) 
      -- 	branch_block_stmt_2042/bb_14_bbx_xnph7x_xix_xix_xi33_PhiReq/phi_stmt_2370/$exit
      -- 	branch_block_stmt_2042/bb_14_bbx_xnph7x_xix_xix_xi33_PhiReq/phi_stmt_2370/phi_stmt_2370_sources/$exit
      -- 	branch_block_stmt_2042/bb_14_bbx_xnph7x_xix_xix_xi33_PhiReq/phi_stmt_2370/phi_stmt_2370_req
      -- 
    cp_element_group_1418: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1418"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1411) & cp_elements(1417);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1418), clk => clk, reset => reset); --
    end block;
    phi_stmt_2370_req_16291_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1418), ack => phi_stmt_2370_req_1); -- 
    -- CP-element group 1419 fork  transition  bypass 
    -- predecessors 1406 
    -- successors 1420 1421 
    -- members (4) 
      -- 	branch_block_stmt_2042/bb_14_bbx_xnph7x_xix_xix_xi33_PhiReq/phi_stmt_2376/$entry
      -- 	branch_block_stmt_2042/bb_14_bbx_xnph7x_xix_xix_xi33_PhiReq/phi_stmt_2376/phi_stmt_2376_sources/$entry
      -- 	branch_block_stmt_2042/bb_14_bbx_xnph7x_xix_xix_xi33_PhiReq/phi_stmt_2376/phi_stmt_2376_sources/type_cast_2379/$entry
      -- 	branch_block_stmt_2042/bb_14_bbx_xnph7x_xix_xix_xi33_PhiReq/phi_stmt_2376/phi_stmt_2376_sources/type_cast_2379/SplitProtocol/$entry
      -- 
    cp_elements(1419) <= cp_elements(1406);
    -- CP-element group 1420 transition  bypass 
    -- predecessors 1419 
    -- successors 1422 
    -- members (4) 
      -- 	branch_block_stmt_2042/bb_14_bbx_xnph7x_xix_xix_xi33_PhiReq/phi_stmt_2376/phi_stmt_2376_sources/type_cast_2379/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_2042/bb_14_bbx_xnph7x_xix_xix_xi33_PhiReq/phi_stmt_2376/phi_stmt_2376_sources/type_cast_2379/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_2042/bb_14_bbx_xnph7x_xix_xix_xi33_PhiReq/phi_stmt_2376/phi_stmt_2376_sources/type_cast_2379/SplitProtocol/Sample/rr
      -- 	branch_block_stmt_2042/bb_14_bbx_xnph7x_xix_xix_xi33_PhiReq/phi_stmt_2376/phi_stmt_2376_sources/type_cast_2379/SplitProtocol/Sample/ra
      -- 
    cp_elements(1420) <= cp_elements(1419);
    -- CP-element group 1421 transition  bypass 
    -- predecessors 1419 
    -- successors 1422 
    -- members (4) 
      -- 	branch_block_stmt_2042/bb_14_bbx_xnph7x_xix_xix_xi33_PhiReq/phi_stmt_2376/phi_stmt_2376_sources/type_cast_2379/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_2042/bb_14_bbx_xnph7x_xix_xix_xi33_PhiReq/phi_stmt_2376/phi_stmt_2376_sources/type_cast_2379/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_2042/bb_14_bbx_xnph7x_xix_xix_xi33_PhiReq/phi_stmt_2376/phi_stmt_2376_sources/type_cast_2379/SplitProtocol/Update/cr
      -- 	branch_block_stmt_2042/bb_14_bbx_xnph7x_xix_xix_xi33_PhiReq/phi_stmt_2376/phi_stmt_2376_sources/type_cast_2379/SplitProtocol/Update/ca
      -- 
    cp_elements(1421) <= cp_elements(1419);
    -- CP-element group 1422 join  transition  output  bypass 
    -- predecessors 1420 1421 
    -- successors 1423 
    -- members (5) 
      -- 	branch_block_stmt_2042/bb_14_bbx_xnph7x_xix_xix_xi33_PhiReq/phi_stmt_2376/$exit
      -- 	branch_block_stmt_2042/bb_14_bbx_xnph7x_xix_xix_xi33_PhiReq/phi_stmt_2376/phi_stmt_2376_sources/$exit
      -- 	branch_block_stmt_2042/bb_14_bbx_xnph7x_xix_xix_xi33_PhiReq/phi_stmt_2376/phi_stmt_2376_sources/type_cast_2379/$exit
      -- 	branch_block_stmt_2042/bb_14_bbx_xnph7x_xix_xix_xi33_PhiReq/phi_stmt_2376/phi_stmt_2376_sources/type_cast_2379/SplitProtocol/$exit
      -- 	branch_block_stmt_2042/bb_14_bbx_xnph7x_xix_xix_xi33_PhiReq/phi_stmt_2376/phi_stmt_2376_req
      -- 
    cp_element_group_1422: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1422"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1420) & cp_elements(1421);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1422), clk => clk, reset => reset); --
    end block;
    phi_stmt_2376_req_16314_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1422), ack => phi_stmt_2376_req_1); -- 
    -- CP-element group 1423 join  transition  bypass 
    -- predecessors 1418 1422 
    -- successors 1444 
    -- members (1) 
      -- 	branch_block_stmt_2042/bb_14_bbx_xnph7x_xix_xix_xi33_PhiReq/$exit
      -- 
    cp_element_group_1423: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1423"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1418) & cp_elements(1422);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1423), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1424 fork  transition  bypass 
    -- predecessors 351 
    -- successors 1425 1437 
    -- members (1) 
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi39_bbx_xnph7x_xix_xix_xi33_PhiReq/$entry
      -- 
    cp_elements(1424) <= cp_elements(351);
    -- CP-element group 1425 fork  transition  bypass 
    -- predecessors 1424 
    -- successors 1426 1432 
    -- members (2) 
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi39_bbx_xnph7x_xix_xix_xi33_PhiReq/phi_stmt_2370/$entry
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi39_bbx_xnph7x_xix_xix_xi33_PhiReq/phi_stmt_2370/phi_stmt_2370_sources/$entry
      -- 
    cp_elements(1425) <= cp_elements(1424);
    -- CP-element group 1426 fork  transition  bypass 
    -- predecessors 1425 
    -- successors 1427 1429 
    -- members (2) 
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi39_bbx_xnph7x_xix_xix_xi33_PhiReq/phi_stmt_2370/phi_stmt_2370_sources/type_cast_2373/$entry
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi39_bbx_xnph7x_xix_xix_xi33_PhiReq/phi_stmt_2370/phi_stmt_2370_sources/type_cast_2373/SplitProtocol/$entry
      -- 
    cp_elements(1426) <= cp_elements(1425);
    -- CP-element group 1427 transition  output  bypass 
    -- predecessors 1426 
    -- successors 1428 
    -- members (2) 
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi39_bbx_xnph7x_xix_xix_xi33_PhiReq/phi_stmt_2370/phi_stmt_2370_sources/type_cast_2373/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi39_bbx_xnph7x_xix_xix_xi33_PhiReq/phi_stmt_2370/phi_stmt_2370_sources/type_cast_2373/SplitProtocol/Sample/rr
      -- 
    cp_elements(1427) <= cp_elements(1426);
    rr_16333_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1427), ack => type_cast_2373_inst_req_0); -- 
    -- CP-element group 1428 transition  input  bypass 
    -- predecessors 1427 
    -- successors 1431 
    -- members (2) 
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi39_bbx_xnph7x_xix_xix_xi33_PhiReq/phi_stmt_2370/phi_stmt_2370_sources/type_cast_2373/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi39_bbx_xnph7x_xix_xix_xi33_PhiReq/phi_stmt_2370/phi_stmt_2370_sources/type_cast_2373/SplitProtocol/Sample/ra
      -- 
    ra_16334_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2373_inst_ack_0, ack => cp_elements(1428)); -- 
    -- CP-element group 1429 transition  output  bypass 
    -- predecessors 1426 
    -- successors 1430 
    -- members (2) 
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi39_bbx_xnph7x_xix_xix_xi33_PhiReq/phi_stmt_2370/phi_stmt_2370_sources/type_cast_2373/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi39_bbx_xnph7x_xix_xix_xi33_PhiReq/phi_stmt_2370/phi_stmt_2370_sources/type_cast_2373/SplitProtocol/Update/cr
      -- 
    cp_elements(1429) <= cp_elements(1426);
    cr_16338_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1429), ack => type_cast_2373_inst_req_1); -- 
    -- CP-element group 1430 transition  input  bypass 
    -- predecessors 1429 
    -- successors 1431 
    -- members (2) 
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi39_bbx_xnph7x_xix_xix_xi33_PhiReq/phi_stmt_2370/phi_stmt_2370_sources/type_cast_2373/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi39_bbx_xnph7x_xix_xix_xi33_PhiReq/phi_stmt_2370/phi_stmt_2370_sources/type_cast_2373/SplitProtocol/Update/ca
      -- 
    ca_16339_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2373_inst_ack_1, ack => cp_elements(1430)); -- 
    -- CP-element group 1431 join  transition  bypass 
    -- predecessors 1428 1430 
    -- successors 1436 
    -- members (2) 
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi39_bbx_xnph7x_xix_xix_xi33_PhiReq/phi_stmt_2370/phi_stmt_2370_sources/type_cast_2373/$exit
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi39_bbx_xnph7x_xix_xix_xi33_PhiReq/phi_stmt_2370/phi_stmt_2370_sources/type_cast_2373/SplitProtocol/$exit
      -- 
    cp_element_group_1431: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1431"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1428) & cp_elements(1430);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1431), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1432 fork  transition  bypass 
    -- predecessors 1425 
    -- successors 1433 1434 
    -- members (2) 
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi39_bbx_xnph7x_xix_xix_xi33_PhiReq/phi_stmt_2370/phi_stmt_2370_sources/type_cast_2375/$entry
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi39_bbx_xnph7x_xix_xix_xi33_PhiReq/phi_stmt_2370/phi_stmt_2370_sources/type_cast_2375/SplitProtocol/$entry
      -- 
    cp_elements(1432) <= cp_elements(1425);
    -- CP-element group 1433 transition  bypass 
    -- predecessors 1432 
    -- successors 1435 
    -- members (4) 
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi39_bbx_xnph7x_xix_xix_xi33_PhiReq/phi_stmt_2370/phi_stmt_2370_sources/type_cast_2375/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi39_bbx_xnph7x_xix_xix_xi33_PhiReq/phi_stmt_2370/phi_stmt_2370_sources/type_cast_2375/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi39_bbx_xnph7x_xix_xix_xi33_PhiReq/phi_stmt_2370/phi_stmt_2370_sources/type_cast_2375/SplitProtocol/Sample/rr
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi39_bbx_xnph7x_xix_xix_xi33_PhiReq/phi_stmt_2370/phi_stmt_2370_sources/type_cast_2375/SplitProtocol/Sample/ra
      -- 
    cp_elements(1433) <= cp_elements(1432);
    -- CP-element group 1434 transition  bypass 
    -- predecessors 1432 
    -- successors 1435 
    -- members (4) 
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi39_bbx_xnph7x_xix_xix_xi33_PhiReq/phi_stmt_2370/phi_stmt_2370_sources/type_cast_2375/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi39_bbx_xnph7x_xix_xix_xi33_PhiReq/phi_stmt_2370/phi_stmt_2370_sources/type_cast_2375/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi39_bbx_xnph7x_xix_xix_xi33_PhiReq/phi_stmt_2370/phi_stmt_2370_sources/type_cast_2375/SplitProtocol/Update/cr
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi39_bbx_xnph7x_xix_xix_xi33_PhiReq/phi_stmt_2370/phi_stmt_2370_sources/type_cast_2375/SplitProtocol/Update/ca
      -- 
    cp_elements(1434) <= cp_elements(1432);
    -- CP-element group 1435 join  transition  bypass 
    -- predecessors 1433 1434 
    -- successors 1436 
    -- members (2) 
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi39_bbx_xnph7x_xix_xix_xi33_PhiReq/phi_stmt_2370/phi_stmt_2370_sources/type_cast_2375/$exit
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi39_bbx_xnph7x_xix_xix_xi33_PhiReq/phi_stmt_2370/phi_stmt_2370_sources/type_cast_2375/SplitProtocol/$exit
      -- 
    cp_element_group_1435: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1435"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1433) & cp_elements(1434);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1435), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1436 join  transition  output  bypass 
    -- predecessors 1431 1435 
    -- successors 1443 
    -- members (3) 
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi39_bbx_xnph7x_xix_xix_xi33_PhiReq/phi_stmt_2370/$exit
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi39_bbx_xnph7x_xix_xix_xi33_PhiReq/phi_stmt_2370/phi_stmt_2370_sources/$exit
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi39_bbx_xnph7x_xix_xix_xi33_PhiReq/phi_stmt_2370/phi_stmt_2370_req
      -- 
    cp_element_group_1436: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1436"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1431) & cp_elements(1435);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1436), clk => clk, reset => reset); --
    end block;
    phi_stmt_2370_req_16356_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1436), ack => phi_stmt_2370_req_0); -- 
    -- CP-element group 1437 fork  transition  bypass 
    -- predecessors 1424 
    -- successors 1438 1440 
    -- members (4) 
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi39_bbx_xnph7x_xix_xix_xi33_PhiReq/phi_stmt_2376/$entry
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi39_bbx_xnph7x_xix_xix_xi33_PhiReq/phi_stmt_2376/phi_stmt_2376_sources/$entry
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi39_bbx_xnph7x_xix_xix_xi33_PhiReq/phi_stmt_2376/phi_stmt_2376_sources/type_cast_2379/$entry
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi39_bbx_xnph7x_xix_xix_xi33_PhiReq/phi_stmt_2376/phi_stmt_2376_sources/type_cast_2379/SplitProtocol/$entry
      -- 
    cp_elements(1437) <= cp_elements(1424);
    -- CP-element group 1438 transition  output  bypass 
    -- predecessors 1437 
    -- successors 1439 
    -- members (2) 
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi39_bbx_xnph7x_xix_xix_xi33_PhiReq/phi_stmt_2376/phi_stmt_2376_sources/type_cast_2379/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi39_bbx_xnph7x_xix_xix_xi33_PhiReq/phi_stmt_2376/phi_stmt_2376_sources/type_cast_2379/SplitProtocol/Sample/rr
      -- 
    cp_elements(1438) <= cp_elements(1437);
    rr_16372_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1438), ack => type_cast_2379_inst_req_0); -- 
    -- CP-element group 1439 transition  input  bypass 
    -- predecessors 1438 
    -- successors 1442 
    -- members (2) 
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi39_bbx_xnph7x_xix_xix_xi33_PhiReq/phi_stmt_2376/phi_stmt_2376_sources/type_cast_2379/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi39_bbx_xnph7x_xix_xix_xi33_PhiReq/phi_stmt_2376/phi_stmt_2376_sources/type_cast_2379/SplitProtocol/Sample/ra
      -- 
    ra_16373_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2379_inst_ack_0, ack => cp_elements(1439)); -- 
    -- CP-element group 1440 transition  output  bypass 
    -- predecessors 1437 
    -- successors 1441 
    -- members (2) 
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi39_bbx_xnph7x_xix_xix_xi33_PhiReq/phi_stmt_2376/phi_stmt_2376_sources/type_cast_2379/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi39_bbx_xnph7x_xix_xix_xi33_PhiReq/phi_stmt_2376/phi_stmt_2376_sources/type_cast_2379/SplitProtocol/Update/cr
      -- 
    cp_elements(1440) <= cp_elements(1437);
    cr_16377_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1440), ack => type_cast_2379_inst_req_1); -- 
    -- CP-element group 1441 transition  input  bypass 
    -- predecessors 1440 
    -- successors 1442 
    -- members (2) 
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi39_bbx_xnph7x_xix_xix_xi33_PhiReq/phi_stmt_2376/phi_stmt_2376_sources/type_cast_2379/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi39_bbx_xnph7x_xix_xix_xi33_PhiReq/phi_stmt_2376/phi_stmt_2376_sources/type_cast_2379/SplitProtocol/Update/ca
      -- 
    ca_16378_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2379_inst_ack_1, ack => cp_elements(1441)); -- 
    -- CP-element group 1442 join  transition  output  bypass 
    -- predecessors 1439 1441 
    -- successors 1443 
    -- members (5) 
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi39_bbx_xnph7x_xix_xix_xi33_PhiReq/phi_stmt_2376/$exit
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi39_bbx_xnph7x_xix_xix_xi33_PhiReq/phi_stmt_2376/phi_stmt_2376_sources/$exit
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi39_bbx_xnph7x_xix_xix_xi33_PhiReq/phi_stmt_2376/phi_stmt_2376_sources/type_cast_2379/$exit
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi39_bbx_xnph7x_xix_xix_xi33_PhiReq/phi_stmt_2376/phi_stmt_2376_sources/type_cast_2379/SplitProtocol/$exit
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi39_bbx_xnph7x_xix_xix_xi33_PhiReq/phi_stmt_2376/phi_stmt_2376_req
      -- 
    cp_element_group_1442: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1442"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1439) & cp_elements(1441);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1442), clk => clk, reset => reset); --
    end block;
    phi_stmt_2376_req_16379_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1442), ack => phi_stmt_2376_req_0); -- 
    -- CP-element group 1443 join  transition  bypass 
    -- predecessors 1436 1442 
    -- successors 1444 
    -- members (1) 
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi39_bbx_xnph7x_xix_xix_xi33_PhiReq/$exit
      -- 
    cp_element_group_1443: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1443"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1436) & cp_elements(1442);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1443), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1444 merge  place  bypass 
    -- predecessors 1423 1443 
    -- successors 1445 
    -- members (1) 
      -- 	branch_block_stmt_2042/merge_stmt_2369_PhiReqMerge
      -- 
    cp_elements(1444) <= OrReduce(cp_elements(1423) & cp_elements(1443));
    -- CP-element group 1445 fork  transition  bypass 
    -- predecessors 1444 
    -- successors 1446 1447 
    -- members (1) 
      -- 	branch_block_stmt_2042/merge_stmt_2369_PhiAck/$entry
      -- 
    cp_elements(1445) <= cp_elements(1444);
    -- CP-element group 1446 transition  input  bypass 
    -- predecessors 1445 
    -- successors 1448 
    -- members (1) 
      -- 	branch_block_stmt_2042/merge_stmt_2369_PhiAck/phi_stmt_2370_ack
      -- 
    phi_stmt_2370_ack_16384_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2370_ack_0, ack => cp_elements(1446)); -- 
    -- CP-element group 1447 transition  input  bypass 
    -- predecessors 1445 
    -- successors 1448 
    -- members (1) 
      -- 	branch_block_stmt_2042/merge_stmt_2369_PhiAck/phi_stmt_2376_ack
      -- 
    phi_stmt_2376_ack_16385_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2376_ack_0, ack => cp_elements(1447)); -- 
    -- CP-element group 1448 join  transition  bypass 
    -- predecessors 1446 1447 
    -- successors 12 
    -- members (1) 
      -- 	branch_block_stmt_2042/merge_stmt_2369_PhiAck/$exit
      -- 
    cp_element_group_1448: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1448"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1446) & cp_elements(1447);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1448), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1449 fork  transition  bypass 
    -- predecessors 325 
    -- successors 1450 1456 
    -- members (1) 
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi36_bbx_xnphx_xix_xix_xi36_PhiReq/$entry
      -- 
    cp_elements(1449) <= cp_elements(325);
    -- CP-element group 1450 fork  transition  bypass 
    -- predecessors 1449 
    -- successors 1451 1453 
    -- members (4) 
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi36_bbx_xnphx_xix_xix_xi36_PhiReq/phi_stmt_2405/$entry
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi36_bbx_xnphx_xix_xix_xi36_PhiReq/phi_stmt_2405/phi_stmt_2405_sources/$entry
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi36_bbx_xnphx_xix_xix_xi36_PhiReq/phi_stmt_2405/phi_stmt_2405_sources/type_cast_2408/$entry
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi36_bbx_xnphx_xix_xix_xi36_PhiReq/phi_stmt_2405/phi_stmt_2405_sources/type_cast_2408/SplitProtocol/$entry
      -- 
    cp_elements(1450) <= cp_elements(1449);
    -- CP-element group 1451 transition  output  bypass 
    -- predecessors 1450 
    -- successors 1452 
    -- members (2) 
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi36_bbx_xnphx_xix_xix_xi36_PhiReq/phi_stmt_2405/phi_stmt_2405_sources/type_cast_2408/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi36_bbx_xnphx_xix_xix_xi36_PhiReq/phi_stmt_2405/phi_stmt_2405_sources/type_cast_2408/SplitProtocol/Sample/rr
      -- 
    cp_elements(1451) <= cp_elements(1450);
    rr_16416_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1451), ack => type_cast_2408_inst_req_0); -- 
    -- CP-element group 1452 transition  input  bypass 
    -- predecessors 1451 
    -- successors 1455 
    -- members (2) 
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi36_bbx_xnphx_xix_xix_xi36_PhiReq/phi_stmt_2405/phi_stmt_2405_sources/type_cast_2408/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi36_bbx_xnphx_xix_xix_xi36_PhiReq/phi_stmt_2405/phi_stmt_2405_sources/type_cast_2408/SplitProtocol/Sample/ra
      -- 
    ra_16417_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2408_inst_ack_0, ack => cp_elements(1452)); -- 
    -- CP-element group 1453 transition  output  bypass 
    -- predecessors 1450 
    -- successors 1454 
    -- members (2) 
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi36_bbx_xnphx_xix_xix_xi36_PhiReq/phi_stmt_2405/phi_stmt_2405_sources/type_cast_2408/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi36_bbx_xnphx_xix_xix_xi36_PhiReq/phi_stmt_2405/phi_stmt_2405_sources/type_cast_2408/SplitProtocol/Update/cr
      -- 
    cp_elements(1453) <= cp_elements(1450);
    cr_16421_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1453), ack => type_cast_2408_inst_req_1); -- 
    -- CP-element group 1454 transition  input  bypass 
    -- predecessors 1453 
    -- successors 1455 
    -- members (2) 
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi36_bbx_xnphx_xix_xix_xi36_PhiReq/phi_stmt_2405/phi_stmt_2405_sources/type_cast_2408/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi36_bbx_xnphx_xix_xix_xi36_PhiReq/phi_stmt_2405/phi_stmt_2405_sources/type_cast_2408/SplitProtocol/Update/ca
      -- 
    ca_16422_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2408_inst_ack_1, ack => cp_elements(1454)); -- 
    -- CP-element group 1455 join  transition  output  bypass 
    -- predecessors 1452 1454 
    -- successors 1462 
    -- members (5) 
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi36_bbx_xnphx_xix_xix_xi36_PhiReq/phi_stmt_2405/$exit
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi36_bbx_xnphx_xix_xix_xi36_PhiReq/phi_stmt_2405/phi_stmt_2405_sources/$exit
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi36_bbx_xnphx_xix_xix_xi36_PhiReq/phi_stmt_2405/phi_stmt_2405_sources/type_cast_2408/$exit
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi36_bbx_xnphx_xix_xix_xi36_PhiReq/phi_stmt_2405/phi_stmt_2405_sources/type_cast_2408/SplitProtocol/$exit
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi36_bbx_xnphx_xix_xix_xi36_PhiReq/phi_stmt_2405/phi_stmt_2405_req
      -- 
    cp_element_group_1455: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1455"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1452) & cp_elements(1454);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1455), clk => clk, reset => reset); --
    end block;
    phi_stmt_2405_req_16423_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1455), ack => phi_stmt_2405_req_0); -- 
    -- CP-element group 1456 fork  transition  bypass 
    -- predecessors 1449 
    -- successors 1457 1459 
    -- members (4) 
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi36_bbx_xnphx_xix_xix_xi36_PhiReq/phi_stmt_2412/$entry
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi36_bbx_xnphx_xix_xix_xi36_PhiReq/phi_stmt_2412/phi_stmt_2412_sources/$entry
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi36_bbx_xnphx_xix_xix_xi36_PhiReq/phi_stmt_2412/phi_stmt_2412_sources/type_cast_2415/$entry
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi36_bbx_xnphx_xix_xix_xi36_PhiReq/phi_stmt_2412/phi_stmt_2412_sources/type_cast_2415/SplitProtocol/$entry
      -- 
    cp_elements(1456) <= cp_elements(1449);
    -- CP-element group 1457 transition  output  bypass 
    -- predecessors 1456 
    -- successors 1458 
    -- members (2) 
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi36_bbx_xnphx_xix_xix_xi36_PhiReq/phi_stmt_2412/phi_stmt_2412_sources/type_cast_2415/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi36_bbx_xnphx_xix_xix_xi36_PhiReq/phi_stmt_2412/phi_stmt_2412_sources/type_cast_2415/SplitProtocol/Sample/rr
      -- 
    cp_elements(1457) <= cp_elements(1456);
    rr_16439_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1457), ack => type_cast_2415_inst_req_0); -- 
    -- CP-element group 1458 transition  input  bypass 
    -- predecessors 1457 
    -- successors 1461 
    -- members (2) 
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi36_bbx_xnphx_xix_xix_xi36_PhiReq/phi_stmt_2412/phi_stmt_2412_sources/type_cast_2415/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi36_bbx_xnphx_xix_xix_xi36_PhiReq/phi_stmt_2412/phi_stmt_2412_sources/type_cast_2415/SplitProtocol/Sample/ra
      -- 
    ra_16440_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2415_inst_ack_0, ack => cp_elements(1458)); -- 
    -- CP-element group 1459 transition  output  bypass 
    -- predecessors 1456 
    -- successors 1460 
    -- members (2) 
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi36_bbx_xnphx_xix_xix_xi36_PhiReq/phi_stmt_2412/phi_stmt_2412_sources/type_cast_2415/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi36_bbx_xnphx_xix_xix_xi36_PhiReq/phi_stmt_2412/phi_stmt_2412_sources/type_cast_2415/SplitProtocol/Update/cr
      -- 
    cp_elements(1459) <= cp_elements(1456);
    cr_16444_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1459), ack => type_cast_2415_inst_req_1); -- 
    -- CP-element group 1460 transition  input  bypass 
    -- predecessors 1459 
    -- successors 1461 
    -- members (2) 
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi36_bbx_xnphx_xix_xix_xi36_PhiReq/phi_stmt_2412/phi_stmt_2412_sources/type_cast_2415/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi36_bbx_xnphx_xix_xix_xi36_PhiReq/phi_stmt_2412/phi_stmt_2412_sources/type_cast_2415/SplitProtocol/Update/ca
      -- 
    ca_16445_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2415_inst_ack_1, ack => cp_elements(1460)); -- 
    -- CP-element group 1461 join  transition  output  bypass 
    -- predecessors 1458 1460 
    -- successors 1462 
    -- members (5) 
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi36_bbx_xnphx_xix_xix_xi36_PhiReq/phi_stmt_2412/$exit
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi36_bbx_xnphx_xix_xix_xi36_PhiReq/phi_stmt_2412/phi_stmt_2412_sources/$exit
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi36_bbx_xnphx_xix_xix_xi36_PhiReq/phi_stmt_2412/phi_stmt_2412_sources/type_cast_2415/$exit
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi36_bbx_xnphx_xix_xix_xi36_PhiReq/phi_stmt_2412/phi_stmt_2412_sources/type_cast_2415/SplitProtocol/$exit
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi36_bbx_xnphx_xix_xix_xi36_PhiReq/phi_stmt_2412/phi_stmt_2412_req
      -- 
    cp_element_group_1461: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1461"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1458) & cp_elements(1460);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1461), clk => clk, reset => reset); --
    end block;
    phi_stmt_2412_req_16446_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1461), ack => phi_stmt_2412_req_0); -- 
    -- CP-element group 1462 join  transition  bypass 
    -- predecessors 1455 1461 
    -- successors 1473 
    -- members (1) 
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi36_bbx_xnphx_xix_xix_xi36_PhiReq/$exit
      -- 
    cp_element_group_1462: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1462"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1455) & cp_elements(1461);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1462), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1463 fork  transition  bypass 
    -- predecessors 13 
    -- successors 1464 1468 
    -- members (1) 
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi36x_xpreheader_bbx_xnphx_xix_xix_xi36_PhiReq/$entry
      -- 
    cp_elements(1463) <= cp_elements(13);
    -- CP-element group 1464 fork  transition  bypass 
    -- predecessors 1463 
    -- successors 1465 1466 
    -- members (4) 
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi36x_xpreheader_bbx_xnphx_xix_xix_xi36_PhiReq/phi_stmt_2405/$entry
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi36x_xpreheader_bbx_xnphx_xix_xix_xi36_PhiReq/phi_stmt_2405/phi_stmt_2405_sources/$entry
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi36x_xpreheader_bbx_xnphx_xix_xix_xi36_PhiReq/phi_stmt_2405/phi_stmt_2405_sources/type_cast_2408/$entry
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi36x_xpreheader_bbx_xnphx_xix_xix_xi36_PhiReq/phi_stmt_2405/phi_stmt_2405_sources/type_cast_2408/SplitProtocol/$entry
      -- 
    cp_elements(1464) <= cp_elements(1463);
    -- CP-element group 1465 transition  bypass 
    -- predecessors 1464 
    -- successors 1467 
    -- members (4) 
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi36x_xpreheader_bbx_xnphx_xix_xix_xi36_PhiReq/phi_stmt_2405/phi_stmt_2405_sources/type_cast_2408/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi36x_xpreheader_bbx_xnphx_xix_xix_xi36_PhiReq/phi_stmt_2405/phi_stmt_2405_sources/type_cast_2408/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi36x_xpreheader_bbx_xnphx_xix_xix_xi36_PhiReq/phi_stmt_2405/phi_stmt_2405_sources/type_cast_2408/SplitProtocol/Sample/rr
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi36x_xpreheader_bbx_xnphx_xix_xix_xi36_PhiReq/phi_stmt_2405/phi_stmt_2405_sources/type_cast_2408/SplitProtocol/Sample/ra
      -- 
    cp_elements(1465) <= cp_elements(1464);
    -- CP-element group 1466 transition  bypass 
    -- predecessors 1464 
    -- successors 1467 
    -- members (4) 
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi36x_xpreheader_bbx_xnphx_xix_xix_xi36_PhiReq/phi_stmt_2405/phi_stmt_2405_sources/type_cast_2408/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi36x_xpreheader_bbx_xnphx_xix_xix_xi36_PhiReq/phi_stmt_2405/phi_stmt_2405_sources/type_cast_2408/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi36x_xpreheader_bbx_xnphx_xix_xix_xi36_PhiReq/phi_stmt_2405/phi_stmt_2405_sources/type_cast_2408/SplitProtocol/Update/cr
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi36x_xpreheader_bbx_xnphx_xix_xix_xi36_PhiReq/phi_stmt_2405/phi_stmt_2405_sources/type_cast_2408/SplitProtocol/Update/ca
      -- 
    cp_elements(1466) <= cp_elements(1464);
    -- CP-element group 1467 join  transition  output  bypass 
    -- predecessors 1465 1466 
    -- successors 1472 
    -- members (5) 
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi36x_xpreheader_bbx_xnphx_xix_xix_xi36_PhiReq/phi_stmt_2405/$exit
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi36x_xpreheader_bbx_xnphx_xix_xix_xi36_PhiReq/phi_stmt_2405/phi_stmt_2405_sources/$exit
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi36x_xpreheader_bbx_xnphx_xix_xix_xi36_PhiReq/phi_stmt_2405/phi_stmt_2405_sources/type_cast_2408/$exit
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi36x_xpreheader_bbx_xnphx_xix_xix_xi36_PhiReq/phi_stmt_2405/phi_stmt_2405_sources/type_cast_2408/SplitProtocol/$exit
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi36x_xpreheader_bbx_xnphx_xix_xix_xi36_PhiReq/phi_stmt_2405/phi_stmt_2405_req
      -- 
    cp_element_group_1467: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1467"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1465) & cp_elements(1466);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1467), clk => clk, reset => reset); --
    end block;
    phi_stmt_2405_req_16472_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1467), ack => phi_stmt_2405_req_1); -- 
    -- CP-element group 1468 fork  transition  bypass 
    -- predecessors 1463 
    -- successors 1469 1470 
    -- members (4) 
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi36x_xpreheader_bbx_xnphx_xix_xix_xi36_PhiReq/phi_stmt_2412/$entry
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi36x_xpreheader_bbx_xnphx_xix_xix_xi36_PhiReq/phi_stmt_2412/phi_stmt_2412_sources/$entry
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi36x_xpreheader_bbx_xnphx_xix_xix_xi36_PhiReq/phi_stmt_2412/phi_stmt_2412_sources/type_cast_2415/$entry
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi36x_xpreheader_bbx_xnphx_xix_xix_xi36_PhiReq/phi_stmt_2412/phi_stmt_2412_sources/type_cast_2415/SplitProtocol/$entry
      -- 
    cp_elements(1468) <= cp_elements(1463);
    -- CP-element group 1469 transition  bypass 
    -- predecessors 1468 
    -- successors 1471 
    -- members (4) 
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi36x_xpreheader_bbx_xnphx_xix_xix_xi36_PhiReq/phi_stmt_2412/phi_stmt_2412_sources/type_cast_2415/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi36x_xpreheader_bbx_xnphx_xix_xix_xi36_PhiReq/phi_stmt_2412/phi_stmt_2412_sources/type_cast_2415/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi36x_xpreheader_bbx_xnphx_xix_xix_xi36_PhiReq/phi_stmt_2412/phi_stmt_2412_sources/type_cast_2415/SplitProtocol/Sample/rr
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi36x_xpreheader_bbx_xnphx_xix_xix_xi36_PhiReq/phi_stmt_2412/phi_stmt_2412_sources/type_cast_2415/SplitProtocol/Sample/ra
      -- 
    cp_elements(1469) <= cp_elements(1468);
    -- CP-element group 1470 transition  bypass 
    -- predecessors 1468 
    -- successors 1471 
    -- members (4) 
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi36x_xpreheader_bbx_xnphx_xix_xix_xi36_PhiReq/phi_stmt_2412/phi_stmt_2412_sources/type_cast_2415/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi36x_xpreheader_bbx_xnphx_xix_xix_xi36_PhiReq/phi_stmt_2412/phi_stmt_2412_sources/type_cast_2415/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi36x_xpreheader_bbx_xnphx_xix_xix_xi36_PhiReq/phi_stmt_2412/phi_stmt_2412_sources/type_cast_2415/SplitProtocol/Update/cr
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi36x_xpreheader_bbx_xnphx_xix_xix_xi36_PhiReq/phi_stmt_2412/phi_stmt_2412_sources/type_cast_2415/SplitProtocol/Update/ca
      -- 
    cp_elements(1470) <= cp_elements(1468);
    -- CP-element group 1471 join  transition  output  bypass 
    -- predecessors 1469 1470 
    -- successors 1472 
    -- members (5) 
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi36x_xpreheader_bbx_xnphx_xix_xix_xi36_PhiReq/phi_stmt_2412/$exit
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi36x_xpreheader_bbx_xnphx_xix_xix_xi36_PhiReq/phi_stmt_2412/phi_stmt_2412_sources/$exit
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi36x_xpreheader_bbx_xnphx_xix_xix_xi36_PhiReq/phi_stmt_2412/phi_stmt_2412_sources/type_cast_2415/$exit
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi36x_xpreheader_bbx_xnphx_xix_xix_xi36_PhiReq/phi_stmt_2412/phi_stmt_2412_sources/type_cast_2415/SplitProtocol/$exit
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi36x_xpreheader_bbx_xnphx_xix_xix_xi36_PhiReq/phi_stmt_2412/phi_stmt_2412_req
      -- 
    cp_element_group_1471: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1471"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1469) & cp_elements(1470);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1471), clk => clk, reset => reset); --
    end block;
    phi_stmt_2412_req_16495_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1471), ack => phi_stmt_2412_req_1); -- 
    -- CP-element group 1472 join  transition  bypass 
    -- predecessors 1467 1471 
    -- successors 1473 
    -- members (1) 
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi36x_xpreheader_bbx_xnphx_xix_xix_xi36_PhiReq/$exit
      -- 
    cp_element_group_1472: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1472"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1467) & cp_elements(1471);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1472), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1473 merge  place  bypass 
    -- predecessors 1462 1472 
    -- successors 1474 
    -- members (1) 
      -- 	branch_block_stmt_2042/merge_stmt_2404_PhiReqMerge
      -- 
    cp_elements(1473) <= OrReduce(cp_elements(1462) & cp_elements(1472));
    -- CP-element group 1474 fork  transition  bypass 
    -- predecessors 1473 
    -- successors 1475 1476 
    -- members (1) 
      -- 	branch_block_stmt_2042/merge_stmt_2404_PhiAck/$entry
      -- 
    cp_elements(1474) <= cp_elements(1473);
    -- CP-element group 1475 transition  input  bypass 
    -- predecessors 1474 
    -- successors 1477 
    -- members (1) 
      -- 	branch_block_stmt_2042/merge_stmt_2404_PhiAck/phi_stmt_2405_ack
      -- 
    phi_stmt_2405_ack_16500_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2405_ack_0, ack => cp_elements(1475)); -- 
    -- CP-element group 1476 transition  input  bypass 
    -- predecessors 1474 
    -- successors 1477 
    -- members (1) 
      -- 	branch_block_stmt_2042/merge_stmt_2404_PhiAck/phi_stmt_2412_ack
      -- 
    phi_stmt_2412_ack_16501_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2412_ack_0, ack => cp_elements(1476)); -- 
    -- CP-element group 1477 join  transition  bypass 
    -- predecessors 1475 1476 
    -- successors 14 
    -- members (1) 
      -- 	branch_block_stmt_2042/merge_stmt_2404_PhiAck/$exit
      -- 
    cp_element_group_1477: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1477"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1475) & cp_elements(1476);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1477), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1478 fork  transition  bypass 
    -- predecessors 327 
    -- successors 1479 1485 
    -- members (1) 
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi36_xx_x_crit_edgex_xix_xix_xi39x_xloopexit_PhiReq/$entry
      -- 
    cp_elements(1478) <= cp_elements(327);
    -- CP-element group 1479 fork  transition  bypass 
    -- predecessors 1478 
    -- successors 1480 1482 
    -- members (4) 
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi36_xx_x_crit_edgex_xix_xix_xi39x_xloopexit_PhiReq/phi_stmt_2444/$entry
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi36_xx_x_crit_edgex_xix_xix_xi39x_xloopexit_PhiReq/phi_stmt_2444/phi_stmt_2444_sources/$entry
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi36_xx_x_crit_edgex_xix_xix_xi39x_xloopexit_PhiReq/phi_stmt_2444/phi_stmt_2444_sources/type_cast_2447/$entry
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi36_xx_x_crit_edgex_xix_xix_xi39x_xloopexit_PhiReq/phi_stmt_2444/phi_stmt_2444_sources/type_cast_2447/SplitProtocol/$entry
      -- 
    cp_elements(1479) <= cp_elements(1478);
    -- CP-element group 1480 transition  output  bypass 
    -- predecessors 1479 
    -- successors 1481 
    -- members (2) 
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi36_xx_x_crit_edgex_xix_xix_xi39x_xloopexit_PhiReq/phi_stmt_2444/phi_stmt_2444_sources/type_cast_2447/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi36_xx_x_crit_edgex_xix_xix_xi39x_xloopexit_PhiReq/phi_stmt_2444/phi_stmt_2444_sources/type_cast_2447/SplitProtocol/Sample/rr
      -- 
    cp_elements(1480) <= cp_elements(1479);
    rr_16524_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1480), ack => type_cast_2447_inst_req_0); -- 
    -- CP-element group 1481 transition  input  bypass 
    -- predecessors 1480 
    -- successors 1484 
    -- members (2) 
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi36_xx_x_crit_edgex_xix_xix_xi39x_xloopexit_PhiReq/phi_stmt_2444/phi_stmt_2444_sources/type_cast_2447/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi36_xx_x_crit_edgex_xix_xix_xi39x_xloopexit_PhiReq/phi_stmt_2444/phi_stmt_2444_sources/type_cast_2447/SplitProtocol/Sample/ra
      -- 
    ra_16525_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2447_inst_ack_0, ack => cp_elements(1481)); -- 
    -- CP-element group 1482 transition  output  bypass 
    -- predecessors 1479 
    -- successors 1483 
    -- members (2) 
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi36_xx_x_crit_edgex_xix_xix_xi39x_xloopexit_PhiReq/phi_stmt_2444/phi_stmt_2444_sources/type_cast_2447/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi36_xx_x_crit_edgex_xix_xix_xi39x_xloopexit_PhiReq/phi_stmt_2444/phi_stmt_2444_sources/type_cast_2447/SplitProtocol/Update/cr
      -- 
    cp_elements(1482) <= cp_elements(1479);
    cr_16529_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1482), ack => type_cast_2447_inst_req_1); -- 
    -- CP-element group 1483 transition  input  bypass 
    -- predecessors 1482 
    -- successors 1484 
    -- members (2) 
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi36_xx_x_crit_edgex_xix_xix_xi39x_xloopexit_PhiReq/phi_stmt_2444/phi_stmt_2444_sources/type_cast_2447/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi36_xx_x_crit_edgex_xix_xix_xi39x_xloopexit_PhiReq/phi_stmt_2444/phi_stmt_2444_sources/type_cast_2447/SplitProtocol/Update/ca
      -- 
    ca_16530_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2447_inst_ack_1, ack => cp_elements(1483)); -- 
    -- CP-element group 1484 join  transition  output  bypass 
    -- predecessors 1481 1483 
    -- successors 1491 
    -- members (5) 
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi36_xx_x_crit_edgex_xix_xix_xi39x_xloopexit_PhiReq/phi_stmt_2444/$exit
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi36_xx_x_crit_edgex_xix_xix_xi39x_xloopexit_PhiReq/phi_stmt_2444/phi_stmt_2444_sources/$exit
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi36_xx_x_crit_edgex_xix_xix_xi39x_xloopexit_PhiReq/phi_stmt_2444/phi_stmt_2444_sources/type_cast_2447/$exit
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi36_xx_x_crit_edgex_xix_xix_xi39x_xloopexit_PhiReq/phi_stmt_2444/phi_stmt_2444_sources/type_cast_2447/SplitProtocol/$exit
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi36_xx_x_crit_edgex_xix_xix_xi39x_xloopexit_PhiReq/phi_stmt_2444/phi_stmt_2444_req
      -- 
    cp_element_group_1484: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1484"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1481) & cp_elements(1483);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1484), clk => clk, reset => reset); --
    end block;
    phi_stmt_2444_req_16531_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1484), ack => phi_stmt_2444_req_0); -- 
    -- CP-element group 1485 fork  transition  bypass 
    -- predecessors 1478 
    -- successors 1486 1488 
    -- members (4) 
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi36_xx_x_crit_edgex_xix_xix_xi39x_xloopexit_PhiReq/phi_stmt_2448/$entry
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi36_xx_x_crit_edgex_xix_xix_xi39x_xloopexit_PhiReq/phi_stmt_2448/phi_stmt_2448_sources/$entry
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi36_xx_x_crit_edgex_xix_xix_xi39x_xloopexit_PhiReq/phi_stmt_2448/phi_stmt_2448_sources/type_cast_2451/$entry
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi36_xx_x_crit_edgex_xix_xix_xi39x_xloopexit_PhiReq/phi_stmt_2448/phi_stmt_2448_sources/type_cast_2451/SplitProtocol/$entry
      -- 
    cp_elements(1485) <= cp_elements(1478);
    -- CP-element group 1486 transition  output  bypass 
    -- predecessors 1485 
    -- successors 1487 
    -- members (2) 
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi36_xx_x_crit_edgex_xix_xix_xi39x_xloopexit_PhiReq/phi_stmt_2448/phi_stmt_2448_sources/type_cast_2451/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi36_xx_x_crit_edgex_xix_xix_xi39x_xloopexit_PhiReq/phi_stmt_2448/phi_stmt_2448_sources/type_cast_2451/SplitProtocol/Sample/rr
      -- 
    cp_elements(1486) <= cp_elements(1485);
    rr_16547_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1486), ack => type_cast_2451_inst_req_0); -- 
    -- CP-element group 1487 transition  input  bypass 
    -- predecessors 1486 
    -- successors 1490 
    -- members (2) 
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi36_xx_x_crit_edgex_xix_xix_xi39x_xloopexit_PhiReq/phi_stmt_2448/phi_stmt_2448_sources/type_cast_2451/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi36_xx_x_crit_edgex_xix_xix_xi39x_xloopexit_PhiReq/phi_stmt_2448/phi_stmt_2448_sources/type_cast_2451/SplitProtocol/Sample/ra
      -- 
    ra_16548_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2451_inst_ack_0, ack => cp_elements(1487)); -- 
    -- CP-element group 1488 transition  output  bypass 
    -- predecessors 1485 
    -- successors 1489 
    -- members (2) 
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi36_xx_x_crit_edgex_xix_xix_xi39x_xloopexit_PhiReq/phi_stmt_2448/phi_stmt_2448_sources/type_cast_2451/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi36_xx_x_crit_edgex_xix_xix_xi39x_xloopexit_PhiReq/phi_stmt_2448/phi_stmt_2448_sources/type_cast_2451/SplitProtocol/Update/cr
      -- 
    cp_elements(1488) <= cp_elements(1485);
    cr_16552_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1488), ack => type_cast_2451_inst_req_1); -- 
    -- CP-element group 1489 transition  input  bypass 
    -- predecessors 1488 
    -- successors 1490 
    -- members (2) 
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi36_xx_x_crit_edgex_xix_xix_xi39x_xloopexit_PhiReq/phi_stmt_2448/phi_stmt_2448_sources/type_cast_2451/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi36_xx_x_crit_edgex_xix_xix_xi39x_xloopexit_PhiReq/phi_stmt_2448/phi_stmt_2448_sources/type_cast_2451/SplitProtocol/Update/ca
      -- 
    ca_16553_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2451_inst_ack_1, ack => cp_elements(1489)); -- 
    -- CP-element group 1490 join  transition  output  bypass 
    -- predecessors 1487 1489 
    -- successors 1491 
    -- members (5) 
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi36_xx_x_crit_edgex_xix_xix_xi39x_xloopexit_PhiReq/phi_stmt_2448/$exit
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi36_xx_x_crit_edgex_xix_xix_xi39x_xloopexit_PhiReq/phi_stmt_2448/phi_stmt_2448_sources/$exit
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi36_xx_x_crit_edgex_xix_xix_xi39x_xloopexit_PhiReq/phi_stmt_2448/phi_stmt_2448_sources/type_cast_2451/$exit
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi36_xx_x_crit_edgex_xix_xix_xi39x_xloopexit_PhiReq/phi_stmt_2448/phi_stmt_2448_sources/type_cast_2451/SplitProtocol/$exit
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi36_xx_x_crit_edgex_xix_xix_xi39x_xloopexit_PhiReq/phi_stmt_2448/phi_stmt_2448_req
      -- 
    cp_element_group_1490: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1490"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1487) & cp_elements(1489);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1490), clk => clk, reset => reset); --
    end block;
    phi_stmt_2448_req_16554_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1490), ack => phi_stmt_2448_req_0); -- 
    -- CP-element group 1491 join  transition  bypass 
    -- predecessors 1484 1490 
    -- successors 1492 
    -- members (1) 
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi36_xx_x_crit_edgex_xix_xix_xi39x_xloopexit_PhiReq/$exit
      -- 
    cp_element_group_1491: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1491"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1484) & cp_elements(1490);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1491), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1492 place  bypass 
    -- predecessors 1491 
    -- successors 1493 
    -- members (1) 
      -- 	branch_block_stmt_2042/merge_stmt_2443_PhiReqMerge
      -- 
    cp_elements(1492) <= cp_elements(1491);
    -- CP-element group 1493 fork  transition  bypass 
    -- predecessors 1492 
    -- successors 1494 1495 
    -- members (1) 
      -- 	branch_block_stmt_2042/merge_stmt_2443_PhiAck/$entry
      -- 
    cp_elements(1493) <= cp_elements(1492);
    -- CP-element group 1494 transition  input  bypass 
    -- predecessors 1493 
    -- successors 1496 
    -- members (1) 
      -- 	branch_block_stmt_2042/merge_stmt_2443_PhiAck/phi_stmt_2444_ack
      -- 
    phi_stmt_2444_ack_16559_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2444_ack_0, ack => cp_elements(1494)); -- 
    -- CP-element group 1495 transition  input  bypass 
    -- predecessors 1493 
    -- successors 1496 
    -- members (1) 
      -- 	branch_block_stmt_2042/merge_stmt_2443_PhiAck/phi_stmt_2448_ack
      -- 
    phi_stmt_2448_ack_16560_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2448_ack_0, ack => cp_elements(1495)); -- 
    -- CP-element group 1496 join  transition  bypass 
    -- predecessors 1494 1495 
    -- successors 16 
    -- members (1) 
      -- 	branch_block_stmt_2042/merge_stmt_2443_PhiAck/$exit
      -- 
    cp_element_group_1496: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1496"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1494) & cp_elements(1495);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1496), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1497 fork  transition  bypass 
    -- predecessors 305 
    -- successors 1498 1502 
    -- members (1) 
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xix_xi33_xx_x_crit_edgex_xix_xix_xi39_PhiReq/$entry
      -- 
    cp_elements(1497) <= cp_elements(305);
    -- CP-element group 1498 fork  transition  bypass 
    -- predecessors 1497 
    -- successors 1499 1500 
    -- members (4) 
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xix_xi33_xx_x_crit_edgex_xix_xix_xi39_PhiReq/phi_stmt_2455/$entry
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xix_xi33_xx_x_crit_edgex_xix_xix_xi39_PhiReq/phi_stmt_2455/phi_stmt_2455_sources/$entry
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xix_xi33_xx_x_crit_edgex_xix_xix_xi39_PhiReq/phi_stmt_2455/phi_stmt_2455_sources/type_cast_2461/$entry
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xix_xi33_xx_x_crit_edgex_xix_xix_xi39_PhiReq/phi_stmt_2455/phi_stmt_2455_sources/type_cast_2461/SplitProtocol/$entry
      -- 
    cp_elements(1498) <= cp_elements(1497);
    -- CP-element group 1499 transition  bypass 
    -- predecessors 1498 
    -- successors 1501 
    -- members (4) 
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xix_xi33_xx_x_crit_edgex_xix_xix_xi39_PhiReq/phi_stmt_2455/phi_stmt_2455_sources/type_cast_2461/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xix_xi33_xx_x_crit_edgex_xix_xix_xi39_PhiReq/phi_stmt_2455/phi_stmt_2455_sources/type_cast_2461/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xix_xi33_xx_x_crit_edgex_xix_xix_xi39_PhiReq/phi_stmt_2455/phi_stmt_2455_sources/type_cast_2461/SplitProtocol/Sample/rr
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xix_xi33_xx_x_crit_edgex_xix_xix_xi39_PhiReq/phi_stmt_2455/phi_stmt_2455_sources/type_cast_2461/SplitProtocol/Sample/ra
      -- 
    cp_elements(1499) <= cp_elements(1498);
    -- CP-element group 1500 transition  bypass 
    -- predecessors 1498 
    -- successors 1501 
    -- members (4) 
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xix_xi33_xx_x_crit_edgex_xix_xix_xi39_PhiReq/phi_stmt_2455/phi_stmt_2455_sources/type_cast_2461/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xix_xi33_xx_x_crit_edgex_xix_xix_xi39_PhiReq/phi_stmt_2455/phi_stmt_2455_sources/type_cast_2461/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xix_xi33_xx_x_crit_edgex_xix_xix_xi39_PhiReq/phi_stmt_2455/phi_stmt_2455_sources/type_cast_2461/SplitProtocol/Update/cr
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xix_xi33_xx_x_crit_edgex_xix_xix_xi39_PhiReq/phi_stmt_2455/phi_stmt_2455_sources/type_cast_2461/SplitProtocol/Update/ca
      -- 
    cp_elements(1500) <= cp_elements(1498);
    -- CP-element group 1501 join  transition  output  bypass 
    -- predecessors 1499 1500 
    -- successors 1506 
    -- members (5) 
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xix_xi33_xx_x_crit_edgex_xix_xix_xi39_PhiReq/phi_stmt_2455/$exit
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xix_xi33_xx_x_crit_edgex_xix_xix_xi39_PhiReq/phi_stmt_2455/phi_stmt_2455_sources/$exit
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xix_xi33_xx_x_crit_edgex_xix_xix_xi39_PhiReq/phi_stmt_2455/phi_stmt_2455_sources/type_cast_2461/$exit
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xix_xi33_xx_x_crit_edgex_xix_xix_xi39_PhiReq/phi_stmt_2455/phi_stmt_2455_sources/type_cast_2461/SplitProtocol/$exit
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xix_xi33_xx_x_crit_edgex_xix_xix_xi39_PhiReq/phi_stmt_2455/phi_stmt_2455_req
      -- 
    cp_element_group_1501: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1501"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1499) & cp_elements(1500);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1501), clk => clk, reset => reset); --
    end block;
    phi_stmt_2455_req_16586_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1501), ack => phi_stmt_2455_req_0); -- 
    -- CP-element group 1502 fork  transition  bypass 
    -- predecessors 1497 
    -- successors 1503 1504 
    -- members (4) 
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xix_xi33_xx_x_crit_edgex_xix_xix_xi39_PhiReq/phi_stmt_2462/$entry
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xix_xi33_xx_x_crit_edgex_xix_xix_xi39_PhiReq/phi_stmt_2462/phi_stmt_2462_sources/$entry
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xix_xi33_xx_x_crit_edgex_xix_xix_xi39_PhiReq/phi_stmt_2462/phi_stmt_2462_sources/type_cast_2468/$entry
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xix_xi33_xx_x_crit_edgex_xix_xix_xi39_PhiReq/phi_stmt_2462/phi_stmt_2462_sources/type_cast_2468/SplitProtocol/$entry
      -- 
    cp_elements(1502) <= cp_elements(1497);
    -- CP-element group 1503 transition  bypass 
    -- predecessors 1502 
    -- successors 1505 
    -- members (4) 
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xix_xi33_xx_x_crit_edgex_xix_xix_xi39_PhiReq/phi_stmt_2462/phi_stmt_2462_sources/type_cast_2468/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xix_xi33_xx_x_crit_edgex_xix_xix_xi39_PhiReq/phi_stmt_2462/phi_stmt_2462_sources/type_cast_2468/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xix_xi33_xx_x_crit_edgex_xix_xix_xi39_PhiReq/phi_stmt_2462/phi_stmt_2462_sources/type_cast_2468/SplitProtocol/Sample/rr
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xix_xi33_xx_x_crit_edgex_xix_xix_xi39_PhiReq/phi_stmt_2462/phi_stmt_2462_sources/type_cast_2468/SplitProtocol/Sample/ra
      -- 
    cp_elements(1503) <= cp_elements(1502);
    -- CP-element group 1504 transition  bypass 
    -- predecessors 1502 
    -- successors 1505 
    -- members (4) 
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xix_xi33_xx_x_crit_edgex_xix_xix_xi39_PhiReq/phi_stmt_2462/phi_stmt_2462_sources/type_cast_2468/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xix_xi33_xx_x_crit_edgex_xix_xix_xi39_PhiReq/phi_stmt_2462/phi_stmt_2462_sources/type_cast_2468/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xix_xi33_xx_x_crit_edgex_xix_xix_xi39_PhiReq/phi_stmt_2462/phi_stmt_2462_sources/type_cast_2468/SplitProtocol/Update/cr
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xix_xi33_xx_x_crit_edgex_xix_xix_xi39_PhiReq/phi_stmt_2462/phi_stmt_2462_sources/type_cast_2468/SplitProtocol/Update/ca
      -- 
    cp_elements(1504) <= cp_elements(1502);
    -- CP-element group 1505 join  transition  output  bypass 
    -- predecessors 1503 1504 
    -- successors 1506 
    -- members (5) 
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xix_xi33_xx_x_crit_edgex_xix_xix_xi39_PhiReq/phi_stmt_2462/$exit
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xix_xi33_xx_x_crit_edgex_xix_xix_xi39_PhiReq/phi_stmt_2462/phi_stmt_2462_sources/$exit
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xix_xi33_xx_x_crit_edgex_xix_xix_xi39_PhiReq/phi_stmt_2462/phi_stmt_2462_sources/type_cast_2468/$exit
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xix_xi33_xx_x_crit_edgex_xix_xix_xi39_PhiReq/phi_stmt_2462/phi_stmt_2462_sources/type_cast_2468/SplitProtocol/$exit
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xix_xi33_xx_x_crit_edgex_xix_xix_xi39_PhiReq/phi_stmt_2462/phi_stmt_2462_req
      -- 
    cp_element_group_1505: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1505"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1503) & cp_elements(1504);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1505), clk => clk, reset => reset); --
    end block;
    phi_stmt_2462_req_16609_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1505), ack => phi_stmt_2462_req_0); -- 
    -- CP-element group 1506 join  transition  bypass 
    -- predecessors 1501 1505 
    -- successors 1521 
    -- members (1) 
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xix_xi33_xx_x_crit_edgex_xix_xix_xi39_PhiReq/$exit
      -- 
    cp_element_group_1506: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1506"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1501) & cp_elements(1505);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1506), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1507 fork  transition  bypass 
    -- predecessors 16 
    -- successors 1508 1514 
    -- members (1) 
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi39x_xloopexit_xx_x_crit_edgex_xix_xix_xi39_PhiReq/$entry
      -- 
    cp_elements(1507) <= cp_elements(16);
    -- CP-element group 1508 fork  transition  bypass 
    -- predecessors 1507 
    -- successors 1509 1511 
    -- members (4) 
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi39x_xloopexit_xx_x_crit_edgex_xix_xix_xi39_PhiReq/phi_stmt_2455/$entry
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi39x_xloopexit_xx_x_crit_edgex_xix_xix_xi39_PhiReq/phi_stmt_2455/phi_stmt_2455_sources/$entry
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi39x_xloopexit_xx_x_crit_edgex_xix_xix_xi39_PhiReq/phi_stmt_2455/phi_stmt_2455_sources/type_cast_2461/$entry
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi39x_xloopexit_xx_x_crit_edgex_xix_xix_xi39_PhiReq/phi_stmt_2455/phi_stmt_2455_sources/type_cast_2461/SplitProtocol/$entry
      -- 
    cp_elements(1508) <= cp_elements(1507);
    -- CP-element group 1509 transition  output  bypass 
    -- predecessors 1508 
    -- successors 1510 
    -- members (2) 
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi39x_xloopexit_xx_x_crit_edgex_xix_xix_xi39_PhiReq/phi_stmt_2455/phi_stmt_2455_sources/type_cast_2461/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi39x_xloopexit_xx_x_crit_edgex_xix_xix_xi39_PhiReq/phi_stmt_2455/phi_stmt_2455_sources/type_cast_2461/SplitProtocol/Sample/rr
      -- 
    cp_elements(1509) <= cp_elements(1508);
    rr_16628_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1509), ack => type_cast_2461_inst_req_0); -- 
    -- CP-element group 1510 transition  input  bypass 
    -- predecessors 1509 
    -- successors 1513 
    -- members (2) 
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi39x_xloopexit_xx_x_crit_edgex_xix_xix_xi39_PhiReq/phi_stmt_2455/phi_stmt_2455_sources/type_cast_2461/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi39x_xloopexit_xx_x_crit_edgex_xix_xix_xi39_PhiReq/phi_stmt_2455/phi_stmt_2455_sources/type_cast_2461/SplitProtocol/Sample/ra
      -- 
    ra_16629_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2461_inst_ack_0, ack => cp_elements(1510)); -- 
    -- CP-element group 1511 transition  output  bypass 
    -- predecessors 1508 
    -- successors 1512 
    -- members (2) 
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi39x_xloopexit_xx_x_crit_edgex_xix_xix_xi39_PhiReq/phi_stmt_2455/phi_stmt_2455_sources/type_cast_2461/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi39x_xloopexit_xx_x_crit_edgex_xix_xix_xi39_PhiReq/phi_stmt_2455/phi_stmt_2455_sources/type_cast_2461/SplitProtocol/Update/cr
      -- 
    cp_elements(1511) <= cp_elements(1508);
    cr_16633_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1511), ack => type_cast_2461_inst_req_1); -- 
    -- CP-element group 1512 transition  input  bypass 
    -- predecessors 1511 
    -- successors 1513 
    -- members (2) 
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi39x_xloopexit_xx_x_crit_edgex_xix_xix_xi39_PhiReq/phi_stmt_2455/phi_stmt_2455_sources/type_cast_2461/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi39x_xloopexit_xx_x_crit_edgex_xix_xix_xi39_PhiReq/phi_stmt_2455/phi_stmt_2455_sources/type_cast_2461/SplitProtocol/Update/ca
      -- 
    ca_16634_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2461_inst_ack_1, ack => cp_elements(1512)); -- 
    -- CP-element group 1513 join  transition  output  bypass 
    -- predecessors 1510 1512 
    -- successors 1520 
    -- members (5) 
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi39x_xloopexit_xx_x_crit_edgex_xix_xix_xi39_PhiReq/phi_stmt_2455/$exit
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi39x_xloopexit_xx_x_crit_edgex_xix_xix_xi39_PhiReq/phi_stmt_2455/phi_stmt_2455_sources/$exit
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi39x_xloopexit_xx_x_crit_edgex_xix_xix_xi39_PhiReq/phi_stmt_2455/phi_stmt_2455_sources/type_cast_2461/$exit
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi39x_xloopexit_xx_x_crit_edgex_xix_xix_xi39_PhiReq/phi_stmt_2455/phi_stmt_2455_sources/type_cast_2461/SplitProtocol/$exit
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi39x_xloopexit_xx_x_crit_edgex_xix_xix_xi39_PhiReq/phi_stmt_2455/phi_stmt_2455_req
      -- 
    cp_element_group_1513: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1513"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1510) & cp_elements(1512);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1513), clk => clk, reset => reset); --
    end block;
    phi_stmt_2455_req_16635_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1513), ack => phi_stmt_2455_req_1); -- 
    -- CP-element group 1514 fork  transition  bypass 
    -- predecessors 1507 
    -- successors 1515 1517 
    -- members (4) 
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi39x_xloopexit_xx_x_crit_edgex_xix_xix_xi39_PhiReq/phi_stmt_2462/$entry
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi39x_xloopexit_xx_x_crit_edgex_xix_xix_xi39_PhiReq/phi_stmt_2462/phi_stmt_2462_sources/$entry
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi39x_xloopexit_xx_x_crit_edgex_xix_xix_xi39_PhiReq/phi_stmt_2462/phi_stmt_2462_sources/type_cast_2468/$entry
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi39x_xloopexit_xx_x_crit_edgex_xix_xix_xi39_PhiReq/phi_stmt_2462/phi_stmt_2462_sources/type_cast_2468/SplitProtocol/$entry
      -- 
    cp_elements(1514) <= cp_elements(1507);
    -- CP-element group 1515 transition  output  bypass 
    -- predecessors 1514 
    -- successors 1516 
    -- members (2) 
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi39x_xloopexit_xx_x_crit_edgex_xix_xix_xi39_PhiReq/phi_stmt_2462/phi_stmt_2462_sources/type_cast_2468/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi39x_xloopexit_xx_x_crit_edgex_xix_xix_xi39_PhiReq/phi_stmt_2462/phi_stmt_2462_sources/type_cast_2468/SplitProtocol/Sample/rr
      -- 
    cp_elements(1515) <= cp_elements(1514);
    rr_16651_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1515), ack => type_cast_2468_inst_req_0); -- 
    -- CP-element group 1516 transition  input  bypass 
    -- predecessors 1515 
    -- successors 1519 
    -- members (2) 
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi39x_xloopexit_xx_x_crit_edgex_xix_xix_xi39_PhiReq/phi_stmt_2462/phi_stmt_2462_sources/type_cast_2468/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi39x_xloopexit_xx_x_crit_edgex_xix_xix_xi39_PhiReq/phi_stmt_2462/phi_stmt_2462_sources/type_cast_2468/SplitProtocol/Sample/ra
      -- 
    ra_16652_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2468_inst_ack_0, ack => cp_elements(1516)); -- 
    -- CP-element group 1517 transition  output  bypass 
    -- predecessors 1514 
    -- successors 1518 
    -- members (2) 
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi39x_xloopexit_xx_x_crit_edgex_xix_xix_xi39_PhiReq/phi_stmt_2462/phi_stmt_2462_sources/type_cast_2468/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi39x_xloopexit_xx_x_crit_edgex_xix_xix_xi39_PhiReq/phi_stmt_2462/phi_stmt_2462_sources/type_cast_2468/SplitProtocol/Update/cr
      -- 
    cp_elements(1517) <= cp_elements(1514);
    cr_16656_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1517), ack => type_cast_2468_inst_req_1); -- 
    -- CP-element group 1518 transition  input  bypass 
    -- predecessors 1517 
    -- successors 1519 
    -- members (2) 
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi39x_xloopexit_xx_x_crit_edgex_xix_xix_xi39_PhiReq/phi_stmt_2462/phi_stmt_2462_sources/type_cast_2468/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi39x_xloopexit_xx_x_crit_edgex_xix_xix_xi39_PhiReq/phi_stmt_2462/phi_stmt_2462_sources/type_cast_2468/SplitProtocol/Update/ca
      -- 
    ca_16657_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2468_inst_ack_1, ack => cp_elements(1518)); -- 
    -- CP-element group 1519 join  transition  output  bypass 
    -- predecessors 1516 1518 
    -- successors 1520 
    -- members (5) 
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi39x_xloopexit_xx_x_crit_edgex_xix_xix_xi39_PhiReq/phi_stmt_2462/$exit
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi39x_xloopexit_xx_x_crit_edgex_xix_xix_xi39_PhiReq/phi_stmt_2462/phi_stmt_2462_sources/$exit
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi39x_xloopexit_xx_x_crit_edgex_xix_xix_xi39_PhiReq/phi_stmt_2462/phi_stmt_2462_sources/type_cast_2468/$exit
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi39x_xloopexit_xx_x_crit_edgex_xix_xix_xi39_PhiReq/phi_stmt_2462/phi_stmt_2462_sources/type_cast_2468/SplitProtocol/$exit
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi39x_xloopexit_xx_x_crit_edgex_xix_xix_xi39_PhiReq/phi_stmt_2462/phi_stmt_2462_req
      -- 
    cp_element_group_1519: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1519"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1516) & cp_elements(1518);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1519), clk => clk, reset => reset); --
    end block;
    phi_stmt_2462_req_16658_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1519), ack => phi_stmt_2462_req_1); -- 
    -- CP-element group 1520 join  transition  bypass 
    -- predecessors 1513 1519 
    -- successors 1521 
    -- members (1) 
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi39x_xloopexit_xx_x_crit_edgex_xix_xix_xi39_PhiReq/$exit
      -- 
    cp_element_group_1520: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1520"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1513) & cp_elements(1519);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1520), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1521 merge  place  bypass 
    -- predecessors 1506 1520 
    -- successors 1522 
    -- members (1) 
      -- 	branch_block_stmt_2042/merge_stmt_2454_PhiReqMerge
      -- 
    cp_elements(1521) <= OrReduce(cp_elements(1506) & cp_elements(1520));
    -- CP-element group 1522 fork  transition  bypass 
    -- predecessors 1521 
    -- successors 1523 1524 
    -- members (1) 
      -- 	branch_block_stmt_2042/merge_stmt_2454_PhiAck/$entry
      -- 
    cp_elements(1522) <= cp_elements(1521);
    -- CP-element group 1523 transition  input  bypass 
    -- predecessors 1522 
    -- successors 1525 
    -- members (1) 
      -- 	branch_block_stmt_2042/merge_stmt_2454_PhiAck/phi_stmt_2455_ack
      -- 
    phi_stmt_2455_ack_16663_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2455_ack_0, ack => cp_elements(1523)); -- 
    -- CP-element group 1524 transition  input  bypass 
    -- predecessors 1522 
    -- successors 1525 
    -- members (1) 
      -- 	branch_block_stmt_2042/merge_stmt_2454_PhiAck/phi_stmt_2462_ack
      -- 
    phi_stmt_2462_ack_16664_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2462_ack_0, ack => cp_elements(1524)); -- 
    -- CP-element group 1525 join  transition  bypass 
    -- predecessors 1523 1524 
    -- successors 17 
    -- members (1) 
      -- 	branch_block_stmt_2042/merge_stmt_2454_PhiAck/$exit
      -- 
    cp_element_group_1525: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1525"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1523) & cp_elements(1524);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1525), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1526 transition  output  bypass 
    -- predecessors 349 
    -- successors 1527 
    -- members (2) 
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi39_udiv32x_xexitx_xpreheaderx_xix_xi41_PhiReq/phi_stmt_2493/phi_stmt_2493_sources/type_cast_2496/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi39_udiv32x_xexitx_xpreheaderx_xix_xi41_PhiReq/phi_stmt_2493/phi_stmt_2493_sources/type_cast_2496/SplitProtocol/Sample/rr
      -- 
    cp_elements(1526) <= cp_elements(349);
    rr_16687_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1526), ack => type_cast_2496_inst_req_0); -- 
    -- CP-element group 1527 transition  input  bypass 
    -- predecessors 1526 
    -- successors 1530 
    -- members (2) 
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi39_udiv32x_xexitx_xpreheaderx_xix_xi41_PhiReq/phi_stmt_2493/phi_stmt_2493_sources/type_cast_2496/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi39_udiv32x_xexitx_xpreheaderx_xix_xi41_PhiReq/phi_stmt_2493/phi_stmt_2493_sources/type_cast_2496/SplitProtocol/Sample/ra
      -- 
    ra_16688_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2496_inst_ack_0, ack => cp_elements(1527)); -- 
    -- CP-element group 1528 transition  output  bypass 
    -- predecessors 349 
    -- successors 1529 
    -- members (2) 
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi39_udiv32x_xexitx_xpreheaderx_xix_xi41_PhiReq/phi_stmt_2493/phi_stmt_2493_sources/type_cast_2496/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi39_udiv32x_xexitx_xpreheaderx_xix_xi41_PhiReq/phi_stmt_2493/phi_stmt_2493_sources/type_cast_2496/SplitProtocol/Update/cr
      -- 
    cp_elements(1528) <= cp_elements(349);
    cr_16692_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1528), ack => type_cast_2496_inst_req_1); -- 
    -- CP-element group 1529 transition  input  bypass 
    -- predecessors 1528 
    -- successors 1530 
    -- members (2) 
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi39_udiv32x_xexitx_xpreheaderx_xix_xi41_PhiReq/phi_stmt_2493/phi_stmt_2493_sources/type_cast_2496/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi39_udiv32x_xexitx_xpreheaderx_xix_xi41_PhiReq/phi_stmt_2493/phi_stmt_2493_sources/type_cast_2496/SplitProtocol/Update/ca
      -- 
    ca_16693_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2496_inst_ack_1, ack => cp_elements(1529)); -- 
    -- CP-element group 1530 join  transition  place  output  bypass 
    -- predecessors 1527 1529 
    -- successors 1531 
    -- members (8) 
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi39_udiv32x_xexitx_xpreheaderx_xix_xi41_PhiReq/$exit
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi39_udiv32x_xexitx_xpreheaderx_xix_xi41_PhiReq/phi_stmt_2493/$exit
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi39_udiv32x_xexitx_xpreheaderx_xix_xi41_PhiReq/phi_stmt_2493/phi_stmt_2493_sources/$exit
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi39_udiv32x_xexitx_xpreheaderx_xix_xi41_PhiReq/phi_stmt_2493/phi_stmt_2493_sources/type_cast_2496/$exit
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi39_udiv32x_xexitx_xpreheaderx_xix_xi41_PhiReq/phi_stmt_2493/phi_stmt_2493_sources/type_cast_2496/SplitProtocol/$exit
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi39_udiv32x_xexitx_xpreheaderx_xix_xi41_PhiReq/phi_stmt_2493/phi_stmt_2493_req
      -- 	branch_block_stmt_2042/merge_stmt_2492_PhiReqMerge
      -- 	branch_block_stmt_2042/merge_stmt_2492_PhiAck/$entry
      -- 
    cp_element_group_1530: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1530"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1527) & cp_elements(1529);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1530), clk => clk, reset => reset); --
    end block;
    phi_stmt_2493_req_16694_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1530), ack => phi_stmt_2493_req_0); -- 
    -- CP-element group 1531 transition  input  bypass 
    -- predecessors 1530 
    -- successors 19 
    -- members (2) 
      -- 	branch_block_stmt_2042/merge_stmt_2492_PhiAck/$exit
      -- 	branch_block_stmt_2042/merge_stmt_2492_PhiAck/phi_stmt_2493_ack
      -- 
    phi_stmt_2493_ack_16699_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2493_ack_0, ack => cp_elements(1531)); -- 
    -- CP-element group 1532 fork  transition  bypass 
    -- predecessors 423 
    -- successors 1533 1539 
    -- members (1) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi45_udiv32x_xexitx_xix_xi45_PhiReq/$entry
      -- 
    cp_elements(1532) <= cp_elements(423);
    -- CP-element group 1533 fork  transition  bypass 
    -- predecessors 1532 
    -- successors 1534 1536 
    -- members (4) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi45_udiv32x_xexitx_xix_xi45_PhiReq/phi_stmt_2556/$entry
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi45_udiv32x_xexitx_xix_xi45_PhiReq/phi_stmt_2556/phi_stmt_2556_sources/$entry
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi45_udiv32x_xexitx_xix_xi45_PhiReq/phi_stmt_2556/phi_stmt_2556_sources/type_cast_2559/$entry
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi45_udiv32x_xexitx_xix_xi45_PhiReq/phi_stmt_2556/phi_stmt_2556_sources/type_cast_2559/SplitProtocol/$entry
      -- 
    cp_elements(1533) <= cp_elements(1532);
    -- CP-element group 1534 transition  output  bypass 
    -- predecessors 1533 
    -- successors 1535 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi45_udiv32x_xexitx_xix_xi45_PhiReq/phi_stmt_2556/phi_stmt_2556_sources/type_cast_2559/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi45_udiv32x_xexitx_xix_xi45_PhiReq/phi_stmt_2556/phi_stmt_2556_sources/type_cast_2559/SplitProtocol/Sample/rr
      -- 
    cp_elements(1534) <= cp_elements(1533);
    rr_16730_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1534), ack => type_cast_2559_inst_req_0); -- 
    -- CP-element group 1535 transition  input  bypass 
    -- predecessors 1534 
    -- successors 1538 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi45_udiv32x_xexitx_xix_xi45_PhiReq/phi_stmt_2556/phi_stmt_2556_sources/type_cast_2559/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi45_udiv32x_xexitx_xix_xi45_PhiReq/phi_stmt_2556/phi_stmt_2556_sources/type_cast_2559/SplitProtocol/Sample/ra
      -- 
    ra_16731_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2559_inst_ack_0, ack => cp_elements(1535)); -- 
    -- CP-element group 1536 transition  output  bypass 
    -- predecessors 1533 
    -- successors 1537 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi45_udiv32x_xexitx_xix_xi45_PhiReq/phi_stmt_2556/phi_stmt_2556_sources/type_cast_2559/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi45_udiv32x_xexitx_xix_xi45_PhiReq/phi_stmt_2556/phi_stmt_2556_sources/type_cast_2559/SplitProtocol/Update/cr
      -- 
    cp_elements(1536) <= cp_elements(1533);
    cr_16735_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1536), ack => type_cast_2559_inst_req_1); -- 
    -- CP-element group 1537 transition  input  bypass 
    -- predecessors 1536 
    -- successors 1538 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi45_udiv32x_xexitx_xix_xi45_PhiReq/phi_stmt_2556/phi_stmt_2556_sources/type_cast_2559/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi45_udiv32x_xexitx_xix_xi45_PhiReq/phi_stmt_2556/phi_stmt_2556_sources/type_cast_2559/SplitProtocol/Update/ca
      -- 
    ca_16736_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2559_inst_ack_1, ack => cp_elements(1537)); -- 
    -- CP-element group 1538 join  transition  output  bypass 
    -- predecessors 1535 1537 
    -- successors 1551 
    -- members (5) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi45_udiv32x_xexitx_xix_xi45_PhiReq/phi_stmt_2556/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi45_udiv32x_xexitx_xix_xi45_PhiReq/phi_stmt_2556/phi_stmt_2556_sources/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi45_udiv32x_xexitx_xix_xi45_PhiReq/phi_stmt_2556/phi_stmt_2556_sources/type_cast_2559/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi45_udiv32x_xexitx_xix_xi45_PhiReq/phi_stmt_2556/phi_stmt_2556_sources/type_cast_2559/SplitProtocol/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi45_udiv32x_xexitx_xix_xi45_PhiReq/phi_stmt_2556/phi_stmt_2556_req
      -- 
    cp_element_group_1538: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1538"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1535) & cp_elements(1537);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1538), clk => clk, reset => reset); --
    end block;
    phi_stmt_2556_req_16737_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1538), ack => phi_stmt_2556_req_0); -- 
    -- CP-element group 1539 fork  transition  bypass 
    -- predecessors 1532 
    -- successors 1540 1546 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi45_udiv32x_xexitx_xix_xi45_PhiReq/phi_stmt_2563/$entry
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi45_udiv32x_xexitx_xix_xi45_PhiReq/phi_stmt_2563/phi_stmt_2563_sources/$entry
      -- 
    cp_elements(1539) <= cp_elements(1532);
    -- CP-element group 1540 fork  transition  bypass 
    -- predecessors 1539 
    -- successors 1541 1543 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi45_udiv32x_xexitx_xix_xi45_PhiReq/phi_stmt_2563/phi_stmt_2563_sources/type_cast_2566/$entry
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi45_udiv32x_xexitx_xix_xi45_PhiReq/phi_stmt_2563/phi_stmt_2563_sources/type_cast_2566/SplitProtocol/$entry
      -- 
    cp_elements(1540) <= cp_elements(1539);
    -- CP-element group 1541 transition  output  bypass 
    -- predecessors 1540 
    -- successors 1542 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi45_udiv32x_xexitx_xix_xi45_PhiReq/phi_stmt_2563/phi_stmt_2563_sources/type_cast_2566/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi45_udiv32x_xexitx_xix_xi45_PhiReq/phi_stmt_2563/phi_stmt_2563_sources/type_cast_2566/SplitProtocol/Sample/rr
      -- 
    cp_elements(1541) <= cp_elements(1540);
    rr_16753_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1541), ack => type_cast_2566_inst_req_0); -- 
    -- CP-element group 1542 transition  input  bypass 
    -- predecessors 1541 
    -- successors 1545 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi45_udiv32x_xexitx_xix_xi45_PhiReq/phi_stmt_2563/phi_stmt_2563_sources/type_cast_2566/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi45_udiv32x_xexitx_xix_xi45_PhiReq/phi_stmt_2563/phi_stmt_2563_sources/type_cast_2566/SplitProtocol/Sample/ra
      -- 
    ra_16754_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2566_inst_ack_0, ack => cp_elements(1542)); -- 
    -- CP-element group 1543 transition  output  bypass 
    -- predecessors 1540 
    -- successors 1544 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi45_udiv32x_xexitx_xix_xi45_PhiReq/phi_stmt_2563/phi_stmt_2563_sources/type_cast_2566/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi45_udiv32x_xexitx_xix_xi45_PhiReq/phi_stmt_2563/phi_stmt_2563_sources/type_cast_2566/SplitProtocol/Update/cr
      -- 
    cp_elements(1543) <= cp_elements(1540);
    cr_16758_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1543), ack => type_cast_2566_inst_req_1); -- 
    -- CP-element group 1544 transition  input  bypass 
    -- predecessors 1543 
    -- successors 1545 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi45_udiv32x_xexitx_xix_xi45_PhiReq/phi_stmt_2563/phi_stmt_2563_sources/type_cast_2566/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi45_udiv32x_xexitx_xix_xi45_PhiReq/phi_stmt_2563/phi_stmt_2563_sources/type_cast_2566/SplitProtocol/Update/ca
      -- 
    ca_16759_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2566_inst_ack_1, ack => cp_elements(1544)); -- 
    -- CP-element group 1545 join  transition  bypass 
    -- predecessors 1542 1544 
    -- successors 1550 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi45_udiv32x_xexitx_xix_xi45_PhiReq/phi_stmt_2563/phi_stmt_2563_sources/type_cast_2566/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi45_udiv32x_xexitx_xix_xi45_PhiReq/phi_stmt_2563/phi_stmt_2563_sources/type_cast_2566/SplitProtocol/$exit
      -- 
    cp_element_group_1545: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1545"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1542) & cp_elements(1544);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1545), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1546 fork  transition  bypass 
    -- predecessors 1539 
    -- successors 1547 1548 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi45_udiv32x_xexitx_xix_xi45_PhiReq/phi_stmt_2563/phi_stmt_2563_sources/type_cast_2568/$entry
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi45_udiv32x_xexitx_xix_xi45_PhiReq/phi_stmt_2563/phi_stmt_2563_sources/type_cast_2568/SplitProtocol/$entry
      -- 
    cp_elements(1546) <= cp_elements(1539);
    -- CP-element group 1547 transition  bypass 
    -- predecessors 1546 
    -- successors 1549 
    -- members (4) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi45_udiv32x_xexitx_xix_xi45_PhiReq/phi_stmt_2563/phi_stmt_2563_sources/type_cast_2568/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi45_udiv32x_xexitx_xix_xi45_PhiReq/phi_stmt_2563/phi_stmt_2563_sources/type_cast_2568/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi45_udiv32x_xexitx_xix_xi45_PhiReq/phi_stmt_2563/phi_stmt_2563_sources/type_cast_2568/SplitProtocol/Sample/rr
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi45_udiv32x_xexitx_xix_xi45_PhiReq/phi_stmt_2563/phi_stmt_2563_sources/type_cast_2568/SplitProtocol/Sample/ra
      -- 
    cp_elements(1547) <= cp_elements(1546);
    -- CP-element group 1548 transition  bypass 
    -- predecessors 1546 
    -- successors 1549 
    -- members (4) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi45_udiv32x_xexitx_xix_xi45_PhiReq/phi_stmt_2563/phi_stmt_2563_sources/type_cast_2568/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi45_udiv32x_xexitx_xix_xi45_PhiReq/phi_stmt_2563/phi_stmt_2563_sources/type_cast_2568/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi45_udiv32x_xexitx_xix_xi45_PhiReq/phi_stmt_2563/phi_stmt_2563_sources/type_cast_2568/SplitProtocol/Update/cr
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi45_udiv32x_xexitx_xix_xi45_PhiReq/phi_stmt_2563/phi_stmt_2563_sources/type_cast_2568/SplitProtocol/Update/ca
      -- 
    cp_elements(1548) <= cp_elements(1546);
    -- CP-element group 1549 join  transition  bypass 
    -- predecessors 1547 1548 
    -- successors 1550 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi45_udiv32x_xexitx_xix_xi45_PhiReq/phi_stmt_2563/phi_stmt_2563_sources/type_cast_2568/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi45_udiv32x_xexitx_xix_xi45_PhiReq/phi_stmt_2563/phi_stmt_2563_sources/type_cast_2568/SplitProtocol/$exit
      -- 
    cp_element_group_1549: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1549"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1547) & cp_elements(1548);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1549), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1550 join  transition  output  bypass 
    -- predecessors 1545 1549 
    -- successors 1551 
    -- members (3) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi45_udiv32x_xexitx_xix_xi45_PhiReq/phi_stmt_2563/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi45_udiv32x_xexitx_xix_xi45_PhiReq/phi_stmt_2563/phi_stmt_2563_sources/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi45_udiv32x_xexitx_xix_xi45_PhiReq/phi_stmt_2563/phi_stmt_2563_req
      -- 
    cp_element_group_1550: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1550"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1545) & cp_elements(1549);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1550), clk => clk, reset => reset); --
    end block;
    phi_stmt_2563_req_16776_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1550), ack => phi_stmt_2563_req_0); -- 
    -- CP-element group 1551 join  transition  bypass 
    -- predecessors 1538 1550 
    -- successors 1570 
    -- members (1) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi45_udiv32x_xexitx_xix_xi45_PhiReq/$exit
      -- 
    cp_element_group_1551: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1551"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1538) & cp_elements(1550);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1551), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1552 fork  transition  bypass 
    -- predecessors 21 
    -- successors 1553 1557 
    -- members (1) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi45x_xpreheader_udiv32x_xexitx_xix_xi45_PhiReq/$entry
      -- 
    cp_elements(1552) <= cp_elements(21);
    -- CP-element group 1553 fork  transition  bypass 
    -- predecessors 1552 
    -- successors 1554 1555 
    -- members (4) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi45x_xpreheader_udiv32x_xexitx_xix_xi45_PhiReq/phi_stmt_2556/$entry
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi45x_xpreheader_udiv32x_xexitx_xix_xi45_PhiReq/phi_stmt_2556/phi_stmt_2556_sources/$entry
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi45x_xpreheader_udiv32x_xexitx_xix_xi45_PhiReq/phi_stmt_2556/phi_stmt_2556_sources/type_cast_2559/$entry
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi45x_xpreheader_udiv32x_xexitx_xix_xi45_PhiReq/phi_stmt_2556/phi_stmt_2556_sources/type_cast_2559/SplitProtocol/$entry
      -- 
    cp_elements(1553) <= cp_elements(1552);
    -- CP-element group 1554 transition  bypass 
    -- predecessors 1553 
    -- successors 1556 
    -- members (4) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi45x_xpreheader_udiv32x_xexitx_xix_xi45_PhiReq/phi_stmt_2556/phi_stmt_2556_sources/type_cast_2559/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi45x_xpreheader_udiv32x_xexitx_xix_xi45_PhiReq/phi_stmt_2556/phi_stmt_2556_sources/type_cast_2559/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi45x_xpreheader_udiv32x_xexitx_xix_xi45_PhiReq/phi_stmt_2556/phi_stmt_2556_sources/type_cast_2559/SplitProtocol/Sample/rr
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi45x_xpreheader_udiv32x_xexitx_xix_xi45_PhiReq/phi_stmt_2556/phi_stmt_2556_sources/type_cast_2559/SplitProtocol/Sample/ra
      -- 
    cp_elements(1554) <= cp_elements(1553);
    -- CP-element group 1555 transition  bypass 
    -- predecessors 1553 
    -- successors 1556 
    -- members (4) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi45x_xpreheader_udiv32x_xexitx_xix_xi45_PhiReq/phi_stmt_2556/phi_stmt_2556_sources/type_cast_2559/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi45x_xpreheader_udiv32x_xexitx_xix_xi45_PhiReq/phi_stmt_2556/phi_stmt_2556_sources/type_cast_2559/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi45x_xpreheader_udiv32x_xexitx_xix_xi45_PhiReq/phi_stmt_2556/phi_stmt_2556_sources/type_cast_2559/SplitProtocol/Update/cr
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi45x_xpreheader_udiv32x_xexitx_xix_xi45_PhiReq/phi_stmt_2556/phi_stmt_2556_sources/type_cast_2559/SplitProtocol/Update/ca
      -- 
    cp_elements(1555) <= cp_elements(1553);
    -- CP-element group 1556 join  transition  output  bypass 
    -- predecessors 1554 1555 
    -- successors 1569 
    -- members (5) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi45x_xpreheader_udiv32x_xexitx_xix_xi45_PhiReq/phi_stmt_2556/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi45x_xpreheader_udiv32x_xexitx_xix_xi45_PhiReq/phi_stmt_2556/phi_stmt_2556_sources/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi45x_xpreheader_udiv32x_xexitx_xix_xi45_PhiReq/phi_stmt_2556/phi_stmt_2556_sources/type_cast_2559/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi45x_xpreheader_udiv32x_xexitx_xix_xi45_PhiReq/phi_stmt_2556/phi_stmt_2556_sources/type_cast_2559/SplitProtocol/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi45x_xpreheader_udiv32x_xexitx_xix_xi45_PhiReq/phi_stmt_2556/phi_stmt_2556_req
      -- 
    cp_element_group_1556: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1556"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1554) & cp_elements(1555);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1556), clk => clk, reset => reset); --
    end block;
    phi_stmt_2556_req_16802_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1556), ack => phi_stmt_2556_req_1); -- 
    -- CP-element group 1557 fork  transition  bypass 
    -- predecessors 1552 
    -- successors 1558 1562 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi45x_xpreheader_udiv32x_xexitx_xix_xi45_PhiReq/phi_stmt_2563/$entry
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi45x_xpreheader_udiv32x_xexitx_xix_xi45_PhiReq/phi_stmt_2563/phi_stmt_2563_sources/$entry
      -- 
    cp_elements(1557) <= cp_elements(1552);
    -- CP-element group 1558 fork  transition  bypass 
    -- predecessors 1557 
    -- successors 1559 1560 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi45x_xpreheader_udiv32x_xexitx_xix_xi45_PhiReq/phi_stmt_2563/phi_stmt_2563_sources/type_cast_2566/$entry
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi45x_xpreheader_udiv32x_xexitx_xix_xi45_PhiReq/phi_stmt_2563/phi_stmt_2563_sources/type_cast_2566/SplitProtocol/$entry
      -- 
    cp_elements(1558) <= cp_elements(1557);
    -- CP-element group 1559 transition  bypass 
    -- predecessors 1558 
    -- successors 1561 
    -- members (4) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi45x_xpreheader_udiv32x_xexitx_xix_xi45_PhiReq/phi_stmt_2563/phi_stmt_2563_sources/type_cast_2566/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi45x_xpreheader_udiv32x_xexitx_xix_xi45_PhiReq/phi_stmt_2563/phi_stmt_2563_sources/type_cast_2566/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi45x_xpreheader_udiv32x_xexitx_xix_xi45_PhiReq/phi_stmt_2563/phi_stmt_2563_sources/type_cast_2566/SplitProtocol/Sample/rr
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi45x_xpreheader_udiv32x_xexitx_xix_xi45_PhiReq/phi_stmt_2563/phi_stmt_2563_sources/type_cast_2566/SplitProtocol/Sample/ra
      -- 
    cp_elements(1559) <= cp_elements(1558);
    -- CP-element group 1560 transition  bypass 
    -- predecessors 1558 
    -- successors 1561 
    -- members (4) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi45x_xpreheader_udiv32x_xexitx_xix_xi45_PhiReq/phi_stmt_2563/phi_stmt_2563_sources/type_cast_2566/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi45x_xpreheader_udiv32x_xexitx_xix_xi45_PhiReq/phi_stmt_2563/phi_stmt_2563_sources/type_cast_2566/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi45x_xpreheader_udiv32x_xexitx_xix_xi45_PhiReq/phi_stmt_2563/phi_stmt_2563_sources/type_cast_2566/SplitProtocol/Update/cr
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi45x_xpreheader_udiv32x_xexitx_xix_xi45_PhiReq/phi_stmt_2563/phi_stmt_2563_sources/type_cast_2566/SplitProtocol/Update/ca
      -- 
    cp_elements(1560) <= cp_elements(1558);
    -- CP-element group 1561 join  transition  bypass 
    -- predecessors 1559 1560 
    -- successors 1568 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi45x_xpreheader_udiv32x_xexitx_xix_xi45_PhiReq/phi_stmt_2563/phi_stmt_2563_sources/type_cast_2566/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi45x_xpreheader_udiv32x_xexitx_xix_xi45_PhiReq/phi_stmt_2563/phi_stmt_2563_sources/type_cast_2566/SplitProtocol/$exit
      -- 
    cp_element_group_1561: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1561"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1559) & cp_elements(1560);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1561), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1562 fork  transition  bypass 
    -- predecessors 1557 
    -- successors 1563 1565 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi45x_xpreheader_udiv32x_xexitx_xix_xi45_PhiReq/phi_stmt_2563/phi_stmt_2563_sources/type_cast_2568/$entry
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi45x_xpreheader_udiv32x_xexitx_xix_xi45_PhiReq/phi_stmt_2563/phi_stmt_2563_sources/type_cast_2568/SplitProtocol/$entry
      -- 
    cp_elements(1562) <= cp_elements(1557);
    -- CP-element group 1563 transition  output  bypass 
    -- predecessors 1562 
    -- successors 1564 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi45x_xpreheader_udiv32x_xexitx_xix_xi45_PhiReq/phi_stmt_2563/phi_stmt_2563_sources/type_cast_2568/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi45x_xpreheader_udiv32x_xexitx_xix_xi45_PhiReq/phi_stmt_2563/phi_stmt_2563_sources/type_cast_2568/SplitProtocol/Sample/rr
      -- 
    cp_elements(1563) <= cp_elements(1562);
    rr_16834_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1563), ack => type_cast_2568_inst_req_0); -- 
    -- CP-element group 1564 transition  input  bypass 
    -- predecessors 1563 
    -- successors 1567 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi45x_xpreheader_udiv32x_xexitx_xix_xi45_PhiReq/phi_stmt_2563/phi_stmt_2563_sources/type_cast_2568/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi45x_xpreheader_udiv32x_xexitx_xix_xi45_PhiReq/phi_stmt_2563/phi_stmt_2563_sources/type_cast_2568/SplitProtocol/Sample/ra
      -- 
    ra_16835_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2568_inst_ack_0, ack => cp_elements(1564)); -- 
    -- CP-element group 1565 transition  output  bypass 
    -- predecessors 1562 
    -- successors 1566 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi45x_xpreheader_udiv32x_xexitx_xix_xi45_PhiReq/phi_stmt_2563/phi_stmt_2563_sources/type_cast_2568/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi45x_xpreheader_udiv32x_xexitx_xix_xi45_PhiReq/phi_stmt_2563/phi_stmt_2563_sources/type_cast_2568/SplitProtocol/Update/cr
      -- 
    cp_elements(1565) <= cp_elements(1562);
    cr_16839_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1565), ack => type_cast_2568_inst_req_1); -- 
    -- CP-element group 1566 transition  input  bypass 
    -- predecessors 1565 
    -- successors 1567 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi45x_xpreheader_udiv32x_xexitx_xix_xi45_PhiReq/phi_stmt_2563/phi_stmt_2563_sources/type_cast_2568/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi45x_xpreheader_udiv32x_xexitx_xix_xi45_PhiReq/phi_stmt_2563/phi_stmt_2563_sources/type_cast_2568/SplitProtocol/Update/ca
      -- 
    ca_16840_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2568_inst_ack_1, ack => cp_elements(1566)); -- 
    -- CP-element group 1567 join  transition  bypass 
    -- predecessors 1564 1566 
    -- successors 1568 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi45x_xpreheader_udiv32x_xexitx_xix_xi45_PhiReq/phi_stmt_2563/phi_stmt_2563_sources/type_cast_2568/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi45x_xpreheader_udiv32x_xexitx_xix_xi45_PhiReq/phi_stmt_2563/phi_stmt_2563_sources/type_cast_2568/SplitProtocol/$exit
      -- 
    cp_element_group_1567: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1567"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1564) & cp_elements(1566);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1567), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1568 join  transition  output  bypass 
    -- predecessors 1561 1567 
    -- successors 1569 
    -- members (3) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi45x_xpreheader_udiv32x_xexitx_xix_xi45_PhiReq/phi_stmt_2563/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi45x_xpreheader_udiv32x_xexitx_xix_xi45_PhiReq/phi_stmt_2563/phi_stmt_2563_sources/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi45x_xpreheader_udiv32x_xexitx_xix_xi45_PhiReq/phi_stmt_2563/phi_stmt_2563_req
      -- 
    cp_element_group_1568: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1568"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1561) & cp_elements(1567);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1568), clk => clk, reset => reset); --
    end block;
    phi_stmt_2563_req_16841_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1568), ack => phi_stmt_2563_req_1); -- 
    -- CP-element group 1569 join  transition  bypass 
    -- predecessors 1556 1568 
    -- successors 1570 
    -- members (1) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi45x_xpreheader_udiv32x_xexitx_xix_xi45_PhiReq/$exit
      -- 
    cp_element_group_1569: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1569"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1556) & cp_elements(1568);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1569), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1570 merge  place  bypass 
    -- predecessors 1551 1569 
    -- successors 1571 
    -- members (1) 
      -- 	branch_block_stmt_2042/merge_stmt_2555_PhiReqMerge
      -- 
    cp_elements(1570) <= OrReduce(cp_elements(1551) & cp_elements(1569));
    -- CP-element group 1571 fork  transition  bypass 
    -- predecessors 1570 
    -- successors 1572 1573 
    -- members (1) 
      -- 	branch_block_stmt_2042/merge_stmt_2555_PhiAck/$entry
      -- 
    cp_elements(1571) <= cp_elements(1570);
    -- CP-element group 1572 transition  input  bypass 
    -- predecessors 1571 
    -- successors 1574 
    -- members (1) 
      -- 	branch_block_stmt_2042/merge_stmt_2555_PhiAck/phi_stmt_2556_ack
      -- 
    phi_stmt_2556_ack_16846_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2556_ack_0, ack => cp_elements(1572)); -- 
    -- CP-element group 1573 transition  input  bypass 
    -- predecessors 1571 
    -- successors 1574 
    -- members (1) 
      -- 	branch_block_stmt_2042/merge_stmt_2555_PhiAck/phi_stmt_2563_ack
      -- 
    phi_stmt_2563_ack_16847_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2563_ack_0, ack => cp_elements(1573)); -- 
    -- CP-element group 1574 join  transition  bypass 
    -- predecessors 1572 1573 
    -- successors 22 
    -- members (1) 
      -- 	branch_block_stmt_2042/merge_stmt_2555_PhiAck/$exit
      -- 
    cp_element_group_1574: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1574"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1572) & cp_elements(1573);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1574), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1575 fork  transition  bypass 
    -- predecessors 425 
    -- successors 1576 1582 
    -- members (1) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi45_udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi48_PhiReq/$entry
      -- 
    cp_elements(1575) <= cp_elements(425);
    -- CP-element group 1576 fork  transition  bypass 
    -- predecessors 1575 
    -- successors 1577 1579 
    -- members (4) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi45_udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi48_PhiReq/phi_stmt_2614/$entry
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi45_udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi48_PhiReq/phi_stmt_2614/phi_stmt_2614_sources/$entry
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi45_udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi48_PhiReq/phi_stmt_2614/phi_stmt_2614_sources/type_cast_2617/$entry
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi45_udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi48_PhiReq/phi_stmt_2614/phi_stmt_2614_sources/type_cast_2617/SplitProtocol/$entry
      -- 
    cp_elements(1576) <= cp_elements(1575);
    -- CP-element group 1577 transition  output  bypass 
    -- predecessors 1576 
    -- successors 1578 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi45_udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi48_PhiReq/phi_stmt_2614/phi_stmt_2614_sources/type_cast_2617/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi45_udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi48_PhiReq/phi_stmt_2614/phi_stmt_2614_sources/type_cast_2617/SplitProtocol/Sample/rr
      -- 
    cp_elements(1577) <= cp_elements(1576);
    rr_16870_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1577), ack => type_cast_2617_inst_req_0); -- 
    -- CP-element group 1578 transition  input  bypass 
    -- predecessors 1577 
    -- successors 1581 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi45_udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi48_PhiReq/phi_stmt_2614/phi_stmt_2614_sources/type_cast_2617/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi45_udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi48_PhiReq/phi_stmt_2614/phi_stmt_2614_sources/type_cast_2617/SplitProtocol/Sample/ra
      -- 
    ra_16871_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2617_inst_ack_0, ack => cp_elements(1578)); -- 
    -- CP-element group 1579 transition  output  bypass 
    -- predecessors 1576 
    -- successors 1580 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi45_udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi48_PhiReq/phi_stmt_2614/phi_stmt_2614_sources/type_cast_2617/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi45_udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi48_PhiReq/phi_stmt_2614/phi_stmt_2614_sources/type_cast_2617/SplitProtocol/Update/cr
      -- 
    cp_elements(1579) <= cp_elements(1576);
    cr_16875_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1579), ack => type_cast_2617_inst_req_1); -- 
    -- CP-element group 1580 transition  input  bypass 
    -- predecessors 1579 
    -- successors 1581 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi45_udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi48_PhiReq/phi_stmt_2614/phi_stmt_2614_sources/type_cast_2617/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi45_udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi48_PhiReq/phi_stmt_2614/phi_stmt_2614_sources/type_cast_2617/SplitProtocol/Update/ca
      -- 
    ca_16876_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2617_inst_ack_1, ack => cp_elements(1580)); -- 
    -- CP-element group 1581 join  transition  output  bypass 
    -- predecessors 1578 1580 
    -- successors 1588 
    -- members (5) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi45_udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi48_PhiReq/phi_stmt_2614/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi45_udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi48_PhiReq/phi_stmt_2614/phi_stmt_2614_sources/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi45_udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi48_PhiReq/phi_stmt_2614/phi_stmt_2614_sources/type_cast_2617/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi45_udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi48_PhiReq/phi_stmt_2614/phi_stmt_2614_sources/type_cast_2617/SplitProtocol/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi45_udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi48_PhiReq/phi_stmt_2614/phi_stmt_2614_req
      -- 
    cp_element_group_1581: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1581"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1578) & cp_elements(1580);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1581), clk => clk, reset => reset); --
    end block;
    phi_stmt_2614_req_16877_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1581), ack => phi_stmt_2614_req_0); -- 
    -- CP-element group 1582 fork  transition  bypass 
    -- predecessors 1575 
    -- successors 1583 1585 
    -- members (4) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi45_udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi48_PhiReq/phi_stmt_2618/$entry
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi45_udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi48_PhiReq/phi_stmt_2618/phi_stmt_2618_sources/$entry
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi45_udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi48_PhiReq/phi_stmt_2618/phi_stmt_2618_sources/type_cast_2621/$entry
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi45_udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi48_PhiReq/phi_stmt_2618/phi_stmt_2618_sources/type_cast_2621/SplitProtocol/$entry
      -- 
    cp_elements(1582) <= cp_elements(1575);
    -- CP-element group 1583 transition  output  bypass 
    -- predecessors 1582 
    -- successors 1584 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi45_udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi48_PhiReq/phi_stmt_2618/phi_stmt_2618_sources/type_cast_2621/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi45_udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi48_PhiReq/phi_stmt_2618/phi_stmt_2618_sources/type_cast_2621/SplitProtocol/Sample/rr
      -- 
    cp_elements(1583) <= cp_elements(1582);
    rr_16893_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1583), ack => type_cast_2621_inst_req_0); -- 
    -- CP-element group 1584 transition  input  bypass 
    -- predecessors 1583 
    -- successors 1587 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi45_udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi48_PhiReq/phi_stmt_2618/phi_stmt_2618_sources/type_cast_2621/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi45_udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi48_PhiReq/phi_stmt_2618/phi_stmt_2618_sources/type_cast_2621/SplitProtocol/Sample/ra
      -- 
    ra_16894_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2621_inst_ack_0, ack => cp_elements(1584)); -- 
    -- CP-element group 1585 transition  output  bypass 
    -- predecessors 1582 
    -- successors 1586 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi45_udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi48_PhiReq/phi_stmt_2618/phi_stmt_2618_sources/type_cast_2621/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi45_udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi48_PhiReq/phi_stmt_2618/phi_stmt_2618_sources/type_cast_2621/SplitProtocol/Update/cr
      -- 
    cp_elements(1585) <= cp_elements(1582);
    cr_16898_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1585), ack => type_cast_2621_inst_req_1); -- 
    -- CP-element group 1586 transition  input  bypass 
    -- predecessors 1585 
    -- successors 1587 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi45_udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi48_PhiReq/phi_stmt_2618/phi_stmt_2618_sources/type_cast_2621/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi45_udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi48_PhiReq/phi_stmt_2618/phi_stmt_2618_sources/type_cast_2621/SplitProtocol/Update/ca
      -- 
    ca_16899_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2621_inst_ack_1, ack => cp_elements(1586)); -- 
    -- CP-element group 1587 join  transition  output  bypass 
    -- predecessors 1584 1586 
    -- successors 1588 
    -- members (5) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi45_udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi48_PhiReq/phi_stmt_2618/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi45_udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi48_PhiReq/phi_stmt_2618/phi_stmt_2618_sources/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi45_udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi48_PhiReq/phi_stmt_2618/phi_stmt_2618_sources/type_cast_2621/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi45_udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi48_PhiReq/phi_stmt_2618/phi_stmt_2618_sources/type_cast_2621/SplitProtocol/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi45_udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi48_PhiReq/phi_stmt_2618/phi_stmt_2618_req
      -- 
    cp_element_group_1587: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1587"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1584) & cp_elements(1586);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1587), clk => clk, reset => reset); --
    end block;
    phi_stmt_2618_req_16900_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1587), ack => phi_stmt_2618_req_0); -- 
    -- CP-element group 1588 join  transition  bypass 
    -- predecessors 1581 1587 
    -- successors 1589 
    -- members (1) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi45_udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi48_PhiReq/$exit
      -- 
    cp_element_group_1588: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1588"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1581) & cp_elements(1587);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1588), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1589 place  bypass 
    -- predecessors 1588 
    -- successors 1590 
    -- members (1) 
      -- 	branch_block_stmt_2042/merge_stmt_2613_PhiReqMerge
      -- 
    cp_elements(1589) <= cp_elements(1588);
    -- CP-element group 1590 fork  transition  bypass 
    -- predecessors 1589 
    -- successors 1591 1592 
    -- members (1) 
      -- 	branch_block_stmt_2042/merge_stmt_2613_PhiAck/$entry
      -- 
    cp_elements(1590) <= cp_elements(1589);
    -- CP-element group 1591 transition  input  bypass 
    -- predecessors 1590 
    -- successors 1593 
    -- members (1) 
      -- 	branch_block_stmt_2042/merge_stmt_2613_PhiAck/phi_stmt_2614_ack
      -- 
    phi_stmt_2614_ack_16905_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2614_ack_0, ack => cp_elements(1591)); -- 
    -- CP-element group 1592 transition  input  bypass 
    -- predecessors 1590 
    -- successors 1593 
    -- members (1) 
      -- 	branch_block_stmt_2042/merge_stmt_2613_PhiAck/phi_stmt_2618_ack
      -- 
    phi_stmt_2618_ack_16906_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2618_ack_0, ack => cp_elements(1592)); -- 
    -- CP-element group 1593 join  transition  bypass 
    -- predecessors 1591 1592 
    -- successors 24 
    -- members (1) 
      -- 	branch_block_stmt_2042/merge_stmt_2613_PhiAck/$exit
      -- 
    cp_element_group_1593: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1593"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1591) & cp_elements(1592);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1593), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1594 fork  transition  bypass 
    -- predecessors 391 
    -- successors 1595 1607 
    -- members (1) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xpreheaderx_xix_xi41_xx_xcritedgex_xix_xi52_PhiReq/$entry
      -- 
    cp_elements(1594) <= cp_elements(391);
    -- CP-element group 1595 fork  transition  bypass 
    -- predecessors 1594 
    -- successors 1596 1600 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xpreheaderx_xix_xi41_xx_xcritedgex_xix_xi52_PhiReq/phi_stmt_2636/$entry
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xpreheaderx_xix_xi41_xx_xcritedgex_xix_xi52_PhiReq/phi_stmt_2636/phi_stmt_2636_sources/$entry
      -- 
    cp_elements(1595) <= cp_elements(1594);
    -- CP-element group 1596 fork  transition  bypass 
    -- predecessors 1595 
    -- successors 1597 1598 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xpreheaderx_xix_xi41_xx_xcritedgex_xix_xi52_PhiReq/phi_stmt_2636/phi_stmt_2636_sources/type_cast_2639/$entry
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xpreheaderx_xix_xi41_xx_xcritedgex_xix_xi52_PhiReq/phi_stmt_2636/phi_stmt_2636_sources/type_cast_2639/SplitProtocol/$entry
      -- 
    cp_elements(1596) <= cp_elements(1595);
    -- CP-element group 1597 transition  bypass 
    -- predecessors 1596 
    -- successors 1599 
    -- members (4) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xpreheaderx_xix_xi41_xx_xcritedgex_xix_xi52_PhiReq/phi_stmt_2636/phi_stmt_2636_sources/type_cast_2639/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xpreheaderx_xix_xi41_xx_xcritedgex_xix_xi52_PhiReq/phi_stmt_2636/phi_stmt_2636_sources/type_cast_2639/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xpreheaderx_xix_xi41_xx_xcritedgex_xix_xi52_PhiReq/phi_stmt_2636/phi_stmt_2636_sources/type_cast_2639/SplitProtocol/Sample/rr
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xpreheaderx_xix_xi41_xx_xcritedgex_xix_xi52_PhiReq/phi_stmt_2636/phi_stmt_2636_sources/type_cast_2639/SplitProtocol/Sample/ra
      -- 
    cp_elements(1597) <= cp_elements(1596);
    -- CP-element group 1598 transition  bypass 
    -- predecessors 1596 
    -- successors 1599 
    -- members (4) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xpreheaderx_xix_xi41_xx_xcritedgex_xix_xi52_PhiReq/phi_stmt_2636/phi_stmt_2636_sources/type_cast_2639/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xpreheaderx_xix_xi41_xx_xcritedgex_xix_xi52_PhiReq/phi_stmt_2636/phi_stmt_2636_sources/type_cast_2639/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xpreheaderx_xix_xi41_xx_xcritedgex_xix_xi52_PhiReq/phi_stmt_2636/phi_stmt_2636_sources/type_cast_2639/SplitProtocol/Update/cr
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xpreheaderx_xix_xi41_xx_xcritedgex_xix_xi52_PhiReq/phi_stmt_2636/phi_stmt_2636_sources/type_cast_2639/SplitProtocol/Update/ca
      -- 
    cp_elements(1598) <= cp_elements(1596);
    -- CP-element group 1599 join  transition  bypass 
    -- predecessors 1597 1598 
    -- successors 1606 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xpreheaderx_xix_xi41_xx_xcritedgex_xix_xi52_PhiReq/phi_stmt_2636/phi_stmt_2636_sources/type_cast_2639/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xpreheaderx_xix_xi41_xx_xcritedgex_xix_xi52_PhiReq/phi_stmt_2636/phi_stmt_2636_sources/type_cast_2639/SplitProtocol/$exit
      -- 
    cp_element_group_1599: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1599"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1597) & cp_elements(1598);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1599), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1600 fork  transition  bypass 
    -- predecessors 1595 
    -- successors 1601 1603 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xpreheaderx_xix_xi41_xx_xcritedgex_xix_xi52_PhiReq/phi_stmt_2636/phi_stmt_2636_sources/type_cast_2641/$entry
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xpreheaderx_xix_xi41_xx_xcritedgex_xix_xi52_PhiReq/phi_stmt_2636/phi_stmt_2636_sources/type_cast_2641/SplitProtocol/$entry
      -- 
    cp_elements(1600) <= cp_elements(1595);
    -- CP-element group 1601 transition  output  bypass 
    -- predecessors 1600 
    -- successors 1602 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xpreheaderx_xix_xi41_xx_xcritedgex_xix_xi52_PhiReq/phi_stmt_2636/phi_stmt_2636_sources/type_cast_2641/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xpreheaderx_xix_xi41_xx_xcritedgex_xix_xi52_PhiReq/phi_stmt_2636/phi_stmt_2636_sources/type_cast_2641/SplitProtocol/Sample/rr
      -- 
    cp_elements(1601) <= cp_elements(1600);
    rr_16941_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1601), ack => type_cast_2641_inst_req_0); -- 
    -- CP-element group 1602 transition  input  bypass 
    -- predecessors 1601 
    -- successors 1605 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xpreheaderx_xix_xi41_xx_xcritedgex_xix_xi52_PhiReq/phi_stmt_2636/phi_stmt_2636_sources/type_cast_2641/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xpreheaderx_xix_xi41_xx_xcritedgex_xix_xi52_PhiReq/phi_stmt_2636/phi_stmt_2636_sources/type_cast_2641/SplitProtocol/Sample/ra
      -- 
    ra_16942_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2641_inst_ack_0, ack => cp_elements(1602)); -- 
    -- CP-element group 1603 transition  output  bypass 
    -- predecessors 1600 
    -- successors 1604 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xpreheaderx_xix_xi41_xx_xcritedgex_xix_xi52_PhiReq/phi_stmt_2636/phi_stmt_2636_sources/type_cast_2641/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xpreheaderx_xix_xi41_xx_xcritedgex_xix_xi52_PhiReq/phi_stmt_2636/phi_stmt_2636_sources/type_cast_2641/SplitProtocol/Update/cr
      -- 
    cp_elements(1603) <= cp_elements(1600);
    cr_16946_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1603), ack => type_cast_2641_inst_req_1); -- 
    -- CP-element group 1604 transition  input  bypass 
    -- predecessors 1603 
    -- successors 1605 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xpreheaderx_xix_xi41_xx_xcritedgex_xix_xi52_PhiReq/phi_stmt_2636/phi_stmt_2636_sources/type_cast_2641/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xpreheaderx_xix_xi41_xx_xcritedgex_xix_xi52_PhiReq/phi_stmt_2636/phi_stmt_2636_sources/type_cast_2641/SplitProtocol/Update/ca
      -- 
    ca_16947_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2641_inst_ack_1, ack => cp_elements(1604)); -- 
    -- CP-element group 1605 join  transition  bypass 
    -- predecessors 1602 1604 
    -- successors 1606 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xpreheaderx_xix_xi41_xx_xcritedgex_xix_xi52_PhiReq/phi_stmt_2636/phi_stmt_2636_sources/type_cast_2641/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xpreheaderx_xix_xi41_xx_xcritedgex_xix_xi52_PhiReq/phi_stmt_2636/phi_stmt_2636_sources/type_cast_2641/SplitProtocol/$exit
      -- 
    cp_element_group_1605: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1605"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1602) & cp_elements(1604);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1605), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1606 join  transition  output  bypass 
    -- predecessors 1599 1605 
    -- successors 1619 
    -- members (3) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xpreheaderx_xix_xi41_xx_xcritedgex_xix_xi52_PhiReq/phi_stmt_2636/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xpreheaderx_xix_xi41_xx_xcritedgex_xix_xi52_PhiReq/phi_stmt_2636/phi_stmt_2636_sources/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xpreheaderx_xix_xi41_xx_xcritedgex_xix_xi52_PhiReq/phi_stmt_2636/phi_stmt_2636_req
      -- 
    cp_element_group_1606: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1606"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1599) & cp_elements(1605);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1606), clk => clk, reset => reset); --
    end block;
    phi_stmt_2636_req_16948_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1606), ack => phi_stmt_2636_req_1); -- 
    -- CP-element group 1607 fork  transition  bypass 
    -- predecessors 1594 
    -- successors 1608 1612 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xpreheaderx_xix_xi41_xx_xcritedgex_xix_xi52_PhiReq/phi_stmt_2642/$entry
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xpreheaderx_xix_xi41_xx_xcritedgex_xix_xi52_PhiReq/phi_stmt_2642/phi_stmt_2642_sources/$entry
      -- 
    cp_elements(1607) <= cp_elements(1594);
    -- CP-element group 1608 fork  transition  bypass 
    -- predecessors 1607 
    -- successors 1609 1610 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xpreheaderx_xix_xi41_xx_xcritedgex_xix_xi52_PhiReq/phi_stmt_2642/phi_stmt_2642_sources/type_cast_2645/$entry
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xpreheaderx_xix_xi41_xx_xcritedgex_xix_xi52_PhiReq/phi_stmt_2642/phi_stmt_2642_sources/type_cast_2645/SplitProtocol/$entry
      -- 
    cp_elements(1608) <= cp_elements(1607);
    -- CP-element group 1609 transition  bypass 
    -- predecessors 1608 
    -- successors 1611 
    -- members (4) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xpreheaderx_xix_xi41_xx_xcritedgex_xix_xi52_PhiReq/phi_stmt_2642/phi_stmt_2642_sources/type_cast_2645/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xpreheaderx_xix_xi41_xx_xcritedgex_xix_xi52_PhiReq/phi_stmt_2642/phi_stmt_2642_sources/type_cast_2645/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xpreheaderx_xix_xi41_xx_xcritedgex_xix_xi52_PhiReq/phi_stmt_2642/phi_stmt_2642_sources/type_cast_2645/SplitProtocol/Sample/rr
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xpreheaderx_xix_xi41_xx_xcritedgex_xix_xi52_PhiReq/phi_stmt_2642/phi_stmt_2642_sources/type_cast_2645/SplitProtocol/Sample/ra
      -- 
    cp_elements(1609) <= cp_elements(1608);
    -- CP-element group 1610 transition  bypass 
    -- predecessors 1608 
    -- successors 1611 
    -- members (4) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xpreheaderx_xix_xi41_xx_xcritedgex_xix_xi52_PhiReq/phi_stmt_2642/phi_stmt_2642_sources/type_cast_2645/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xpreheaderx_xix_xi41_xx_xcritedgex_xix_xi52_PhiReq/phi_stmt_2642/phi_stmt_2642_sources/type_cast_2645/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xpreheaderx_xix_xi41_xx_xcritedgex_xix_xi52_PhiReq/phi_stmt_2642/phi_stmt_2642_sources/type_cast_2645/SplitProtocol/Update/cr
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xpreheaderx_xix_xi41_xx_xcritedgex_xix_xi52_PhiReq/phi_stmt_2642/phi_stmt_2642_sources/type_cast_2645/SplitProtocol/Update/ca
      -- 
    cp_elements(1610) <= cp_elements(1608);
    -- CP-element group 1611 join  transition  bypass 
    -- predecessors 1609 1610 
    -- successors 1618 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xpreheaderx_xix_xi41_xx_xcritedgex_xix_xi52_PhiReq/phi_stmt_2642/phi_stmt_2642_sources/type_cast_2645/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xpreheaderx_xix_xi41_xx_xcritedgex_xix_xi52_PhiReq/phi_stmt_2642/phi_stmt_2642_sources/type_cast_2645/SplitProtocol/$exit
      -- 
    cp_element_group_1611: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1611"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1609) & cp_elements(1610);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1611), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1612 fork  transition  bypass 
    -- predecessors 1607 
    -- successors 1613 1615 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xpreheaderx_xix_xi41_xx_xcritedgex_xix_xi52_PhiReq/phi_stmt_2642/phi_stmt_2642_sources/type_cast_2647/$entry
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xpreheaderx_xix_xi41_xx_xcritedgex_xix_xi52_PhiReq/phi_stmt_2642/phi_stmt_2642_sources/type_cast_2647/SplitProtocol/$entry
      -- 
    cp_elements(1612) <= cp_elements(1607);
    -- CP-element group 1613 transition  output  bypass 
    -- predecessors 1612 
    -- successors 1614 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xpreheaderx_xix_xi41_xx_xcritedgex_xix_xi52_PhiReq/phi_stmt_2642/phi_stmt_2642_sources/type_cast_2647/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xpreheaderx_xix_xi41_xx_xcritedgex_xix_xi52_PhiReq/phi_stmt_2642/phi_stmt_2642_sources/type_cast_2647/SplitProtocol/Sample/rr
      -- 
    cp_elements(1613) <= cp_elements(1612);
    rr_16980_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1613), ack => type_cast_2647_inst_req_0); -- 
    -- CP-element group 1614 transition  input  bypass 
    -- predecessors 1613 
    -- successors 1617 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xpreheaderx_xix_xi41_xx_xcritedgex_xix_xi52_PhiReq/phi_stmt_2642/phi_stmt_2642_sources/type_cast_2647/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xpreheaderx_xix_xi41_xx_xcritedgex_xix_xi52_PhiReq/phi_stmt_2642/phi_stmt_2642_sources/type_cast_2647/SplitProtocol/Sample/ra
      -- 
    ra_16981_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2647_inst_ack_0, ack => cp_elements(1614)); -- 
    -- CP-element group 1615 transition  output  bypass 
    -- predecessors 1612 
    -- successors 1616 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xpreheaderx_xix_xi41_xx_xcritedgex_xix_xi52_PhiReq/phi_stmt_2642/phi_stmt_2642_sources/type_cast_2647/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xpreheaderx_xix_xi41_xx_xcritedgex_xix_xi52_PhiReq/phi_stmt_2642/phi_stmt_2642_sources/type_cast_2647/SplitProtocol/Update/cr
      -- 
    cp_elements(1615) <= cp_elements(1612);
    cr_16985_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1615), ack => type_cast_2647_inst_req_1); -- 
    -- CP-element group 1616 transition  input  bypass 
    -- predecessors 1615 
    -- successors 1617 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xpreheaderx_xix_xi41_xx_xcritedgex_xix_xi52_PhiReq/phi_stmt_2642/phi_stmt_2642_sources/type_cast_2647/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xpreheaderx_xix_xi41_xx_xcritedgex_xix_xi52_PhiReq/phi_stmt_2642/phi_stmt_2642_sources/type_cast_2647/SplitProtocol/Update/ca
      -- 
    ca_16986_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2647_inst_ack_1, ack => cp_elements(1616)); -- 
    -- CP-element group 1617 join  transition  bypass 
    -- predecessors 1614 1616 
    -- successors 1618 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xpreheaderx_xix_xi41_xx_xcritedgex_xix_xi52_PhiReq/phi_stmt_2642/phi_stmt_2642_sources/type_cast_2647/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xpreheaderx_xix_xi41_xx_xcritedgex_xix_xi52_PhiReq/phi_stmt_2642/phi_stmt_2642_sources/type_cast_2647/SplitProtocol/$exit
      -- 
    cp_element_group_1617: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1617"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1614) & cp_elements(1616);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1617), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1618 join  transition  output  bypass 
    -- predecessors 1611 1617 
    -- successors 1619 
    -- members (3) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xpreheaderx_xix_xi41_xx_xcritedgex_xix_xi52_PhiReq/phi_stmt_2642/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xpreheaderx_xix_xi41_xx_xcritedgex_xix_xi52_PhiReq/phi_stmt_2642/phi_stmt_2642_sources/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xpreheaderx_xix_xi41_xx_xcritedgex_xix_xi52_PhiReq/phi_stmt_2642/phi_stmt_2642_req
      -- 
    cp_element_group_1618: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1618"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1611) & cp_elements(1617);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1618), clk => clk, reset => reset); --
    end block;
    phi_stmt_2642_req_16987_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1618), ack => phi_stmt_2642_req_1); -- 
    -- CP-element group 1619 join  transition  bypass 
    -- predecessors 1606 1618 
    -- successors 1646 
    -- members (1) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xpreheaderx_xix_xi41_xx_xcritedgex_xix_xi52_PhiReq/$exit
      -- 
    cp_element_group_1619: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1619"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1606) & cp_elements(1618);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1619), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1620 fork  transition  bypass 
    -- predecessors 435 
    -- successors 1621 1633 
    -- members (1) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi48_xx_xcritedgex_xix_xi52_PhiReq/$entry
      -- 
    cp_elements(1620) <= cp_elements(435);
    -- CP-element group 1621 fork  transition  bypass 
    -- predecessors 1620 
    -- successors 1622 1628 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi48_xx_xcritedgex_xix_xi52_PhiReq/phi_stmt_2636/$entry
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi48_xx_xcritedgex_xix_xi52_PhiReq/phi_stmt_2636/phi_stmt_2636_sources/$entry
      -- 
    cp_elements(1621) <= cp_elements(1620);
    -- CP-element group 1622 fork  transition  bypass 
    -- predecessors 1621 
    -- successors 1623 1625 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi48_xx_xcritedgex_xix_xi52_PhiReq/phi_stmt_2636/phi_stmt_2636_sources/type_cast_2639/$entry
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi48_xx_xcritedgex_xix_xi52_PhiReq/phi_stmt_2636/phi_stmt_2636_sources/type_cast_2639/SplitProtocol/$entry
      -- 
    cp_elements(1622) <= cp_elements(1621);
    -- CP-element group 1623 transition  output  bypass 
    -- predecessors 1622 
    -- successors 1624 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi48_xx_xcritedgex_xix_xi52_PhiReq/phi_stmt_2636/phi_stmt_2636_sources/type_cast_2639/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi48_xx_xcritedgex_xix_xi52_PhiReq/phi_stmt_2636/phi_stmt_2636_sources/type_cast_2639/SplitProtocol/Sample/rr
      -- 
    cp_elements(1623) <= cp_elements(1622);
    rr_17006_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1623), ack => type_cast_2639_inst_req_0); -- 
    -- CP-element group 1624 transition  input  bypass 
    -- predecessors 1623 
    -- successors 1627 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi48_xx_xcritedgex_xix_xi52_PhiReq/phi_stmt_2636/phi_stmt_2636_sources/type_cast_2639/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi48_xx_xcritedgex_xix_xi52_PhiReq/phi_stmt_2636/phi_stmt_2636_sources/type_cast_2639/SplitProtocol/Sample/ra
      -- 
    ra_17007_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2639_inst_ack_0, ack => cp_elements(1624)); -- 
    -- CP-element group 1625 transition  output  bypass 
    -- predecessors 1622 
    -- successors 1626 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi48_xx_xcritedgex_xix_xi52_PhiReq/phi_stmt_2636/phi_stmt_2636_sources/type_cast_2639/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi48_xx_xcritedgex_xix_xi52_PhiReq/phi_stmt_2636/phi_stmt_2636_sources/type_cast_2639/SplitProtocol/Update/cr
      -- 
    cp_elements(1625) <= cp_elements(1622);
    cr_17011_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1625), ack => type_cast_2639_inst_req_1); -- 
    -- CP-element group 1626 transition  input  bypass 
    -- predecessors 1625 
    -- successors 1627 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi48_xx_xcritedgex_xix_xi52_PhiReq/phi_stmt_2636/phi_stmt_2636_sources/type_cast_2639/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi48_xx_xcritedgex_xix_xi52_PhiReq/phi_stmt_2636/phi_stmt_2636_sources/type_cast_2639/SplitProtocol/Update/ca
      -- 
    ca_17012_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2639_inst_ack_1, ack => cp_elements(1626)); -- 
    -- CP-element group 1627 join  transition  bypass 
    -- predecessors 1624 1626 
    -- successors 1632 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi48_xx_xcritedgex_xix_xi52_PhiReq/phi_stmt_2636/phi_stmt_2636_sources/type_cast_2639/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi48_xx_xcritedgex_xix_xi52_PhiReq/phi_stmt_2636/phi_stmt_2636_sources/type_cast_2639/SplitProtocol/$exit
      -- 
    cp_element_group_1627: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1627"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1624) & cp_elements(1626);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1627), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1628 fork  transition  bypass 
    -- predecessors 1621 
    -- successors 1629 1630 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi48_xx_xcritedgex_xix_xi52_PhiReq/phi_stmt_2636/phi_stmt_2636_sources/type_cast_2641/$entry
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi48_xx_xcritedgex_xix_xi52_PhiReq/phi_stmt_2636/phi_stmt_2636_sources/type_cast_2641/SplitProtocol/$entry
      -- 
    cp_elements(1628) <= cp_elements(1621);
    -- CP-element group 1629 transition  bypass 
    -- predecessors 1628 
    -- successors 1631 
    -- members (4) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi48_xx_xcritedgex_xix_xi52_PhiReq/phi_stmt_2636/phi_stmt_2636_sources/type_cast_2641/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi48_xx_xcritedgex_xix_xi52_PhiReq/phi_stmt_2636/phi_stmt_2636_sources/type_cast_2641/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi48_xx_xcritedgex_xix_xi52_PhiReq/phi_stmt_2636/phi_stmt_2636_sources/type_cast_2641/SplitProtocol/Sample/rr
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi48_xx_xcritedgex_xix_xi52_PhiReq/phi_stmt_2636/phi_stmt_2636_sources/type_cast_2641/SplitProtocol/Sample/ra
      -- 
    cp_elements(1629) <= cp_elements(1628);
    -- CP-element group 1630 transition  bypass 
    -- predecessors 1628 
    -- successors 1631 
    -- members (4) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi48_xx_xcritedgex_xix_xi52_PhiReq/phi_stmt_2636/phi_stmt_2636_sources/type_cast_2641/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi48_xx_xcritedgex_xix_xi52_PhiReq/phi_stmt_2636/phi_stmt_2636_sources/type_cast_2641/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi48_xx_xcritedgex_xix_xi52_PhiReq/phi_stmt_2636/phi_stmt_2636_sources/type_cast_2641/SplitProtocol/Update/cr
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi48_xx_xcritedgex_xix_xi52_PhiReq/phi_stmt_2636/phi_stmt_2636_sources/type_cast_2641/SplitProtocol/Update/ca
      -- 
    cp_elements(1630) <= cp_elements(1628);
    -- CP-element group 1631 join  transition  bypass 
    -- predecessors 1629 1630 
    -- successors 1632 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi48_xx_xcritedgex_xix_xi52_PhiReq/phi_stmt_2636/phi_stmt_2636_sources/type_cast_2641/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi48_xx_xcritedgex_xix_xi52_PhiReq/phi_stmt_2636/phi_stmt_2636_sources/type_cast_2641/SplitProtocol/$exit
      -- 
    cp_element_group_1631: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1631"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1629) & cp_elements(1630);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1631), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1632 join  transition  output  bypass 
    -- predecessors 1627 1631 
    -- successors 1645 
    -- members (3) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi48_xx_xcritedgex_xix_xi52_PhiReq/phi_stmt_2636/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi48_xx_xcritedgex_xix_xi52_PhiReq/phi_stmt_2636/phi_stmt_2636_sources/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi48_xx_xcritedgex_xix_xi52_PhiReq/phi_stmt_2636/phi_stmt_2636_req
      -- 
    cp_element_group_1632: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1632"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1627) & cp_elements(1631);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1632), clk => clk, reset => reset); --
    end block;
    phi_stmt_2636_req_17029_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1632), ack => phi_stmt_2636_req_0); -- 
    -- CP-element group 1633 fork  transition  bypass 
    -- predecessors 1620 
    -- successors 1634 1640 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi48_xx_xcritedgex_xix_xi52_PhiReq/phi_stmt_2642/$entry
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi48_xx_xcritedgex_xix_xi52_PhiReq/phi_stmt_2642/phi_stmt_2642_sources/$entry
      -- 
    cp_elements(1633) <= cp_elements(1620);
    -- CP-element group 1634 fork  transition  bypass 
    -- predecessors 1633 
    -- successors 1635 1637 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi48_xx_xcritedgex_xix_xi52_PhiReq/phi_stmt_2642/phi_stmt_2642_sources/type_cast_2645/$entry
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi48_xx_xcritedgex_xix_xi52_PhiReq/phi_stmt_2642/phi_stmt_2642_sources/type_cast_2645/SplitProtocol/$entry
      -- 
    cp_elements(1634) <= cp_elements(1633);
    -- CP-element group 1635 transition  output  bypass 
    -- predecessors 1634 
    -- successors 1636 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi48_xx_xcritedgex_xix_xi52_PhiReq/phi_stmt_2642/phi_stmt_2642_sources/type_cast_2645/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi48_xx_xcritedgex_xix_xi52_PhiReq/phi_stmt_2642/phi_stmt_2642_sources/type_cast_2645/SplitProtocol/Sample/rr
      -- 
    cp_elements(1635) <= cp_elements(1634);
    rr_17045_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1635), ack => type_cast_2645_inst_req_0); -- 
    -- CP-element group 1636 transition  input  bypass 
    -- predecessors 1635 
    -- successors 1639 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi48_xx_xcritedgex_xix_xi52_PhiReq/phi_stmt_2642/phi_stmt_2642_sources/type_cast_2645/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi48_xx_xcritedgex_xix_xi52_PhiReq/phi_stmt_2642/phi_stmt_2642_sources/type_cast_2645/SplitProtocol/Sample/ra
      -- 
    ra_17046_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2645_inst_ack_0, ack => cp_elements(1636)); -- 
    -- CP-element group 1637 transition  output  bypass 
    -- predecessors 1634 
    -- successors 1638 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi48_xx_xcritedgex_xix_xi52_PhiReq/phi_stmt_2642/phi_stmt_2642_sources/type_cast_2645/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi48_xx_xcritedgex_xix_xi52_PhiReq/phi_stmt_2642/phi_stmt_2642_sources/type_cast_2645/SplitProtocol/Update/cr
      -- 
    cp_elements(1637) <= cp_elements(1634);
    cr_17050_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1637), ack => type_cast_2645_inst_req_1); -- 
    -- CP-element group 1638 transition  input  bypass 
    -- predecessors 1637 
    -- successors 1639 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi48_xx_xcritedgex_xix_xi52_PhiReq/phi_stmt_2642/phi_stmt_2642_sources/type_cast_2645/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi48_xx_xcritedgex_xix_xi52_PhiReq/phi_stmt_2642/phi_stmt_2642_sources/type_cast_2645/SplitProtocol/Update/ca
      -- 
    ca_17051_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2645_inst_ack_1, ack => cp_elements(1638)); -- 
    -- CP-element group 1639 join  transition  bypass 
    -- predecessors 1636 1638 
    -- successors 1644 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi48_xx_xcritedgex_xix_xi52_PhiReq/phi_stmt_2642/phi_stmt_2642_sources/type_cast_2645/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi48_xx_xcritedgex_xix_xi52_PhiReq/phi_stmt_2642/phi_stmt_2642_sources/type_cast_2645/SplitProtocol/$exit
      -- 
    cp_element_group_1639: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1639"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1636) & cp_elements(1638);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1639), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1640 fork  transition  bypass 
    -- predecessors 1633 
    -- successors 1641 1642 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi48_xx_xcritedgex_xix_xi52_PhiReq/phi_stmt_2642/phi_stmt_2642_sources/type_cast_2647/$entry
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi48_xx_xcritedgex_xix_xi52_PhiReq/phi_stmt_2642/phi_stmt_2642_sources/type_cast_2647/SplitProtocol/$entry
      -- 
    cp_elements(1640) <= cp_elements(1633);
    -- CP-element group 1641 transition  bypass 
    -- predecessors 1640 
    -- successors 1643 
    -- members (4) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi48_xx_xcritedgex_xix_xi52_PhiReq/phi_stmt_2642/phi_stmt_2642_sources/type_cast_2647/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi48_xx_xcritedgex_xix_xi52_PhiReq/phi_stmt_2642/phi_stmt_2642_sources/type_cast_2647/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi48_xx_xcritedgex_xix_xi52_PhiReq/phi_stmt_2642/phi_stmt_2642_sources/type_cast_2647/SplitProtocol/Sample/rr
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi48_xx_xcritedgex_xix_xi52_PhiReq/phi_stmt_2642/phi_stmt_2642_sources/type_cast_2647/SplitProtocol/Sample/ra
      -- 
    cp_elements(1641) <= cp_elements(1640);
    -- CP-element group 1642 transition  bypass 
    -- predecessors 1640 
    -- successors 1643 
    -- members (4) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi48_xx_xcritedgex_xix_xi52_PhiReq/phi_stmt_2642/phi_stmt_2642_sources/type_cast_2647/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi48_xx_xcritedgex_xix_xi52_PhiReq/phi_stmt_2642/phi_stmt_2642_sources/type_cast_2647/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi48_xx_xcritedgex_xix_xi52_PhiReq/phi_stmt_2642/phi_stmt_2642_sources/type_cast_2647/SplitProtocol/Update/cr
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi48_xx_xcritedgex_xix_xi52_PhiReq/phi_stmt_2642/phi_stmt_2642_sources/type_cast_2647/SplitProtocol/Update/ca
      -- 
    cp_elements(1642) <= cp_elements(1640);
    -- CP-element group 1643 join  transition  bypass 
    -- predecessors 1641 1642 
    -- successors 1644 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi48_xx_xcritedgex_xix_xi52_PhiReq/phi_stmt_2642/phi_stmt_2642_sources/type_cast_2647/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi48_xx_xcritedgex_xix_xi52_PhiReq/phi_stmt_2642/phi_stmt_2642_sources/type_cast_2647/SplitProtocol/$exit
      -- 
    cp_element_group_1643: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1643"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1641) & cp_elements(1642);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1643), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1644 join  transition  output  bypass 
    -- predecessors 1639 1643 
    -- successors 1645 
    -- members (3) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi48_xx_xcritedgex_xix_xi52_PhiReq/phi_stmt_2642/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi48_xx_xcritedgex_xix_xi52_PhiReq/phi_stmt_2642/phi_stmt_2642_sources/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi48_xx_xcritedgex_xix_xi52_PhiReq/phi_stmt_2642/phi_stmt_2642_req
      -- 
    cp_element_group_1644: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1644"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1639) & cp_elements(1643);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1644), clk => clk, reset => reset); --
    end block;
    phi_stmt_2642_req_17068_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1644), ack => phi_stmt_2642_req_0); -- 
    -- CP-element group 1645 join  transition  bypass 
    -- predecessors 1632 1644 
    -- successors 1646 
    -- members (1) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi48_xx_xcritedgex_xix_xi52_PhiReq/$exit
      -- 
    cp_element_group_1645: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1645"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1632) & cp_elements(1644);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1645), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1646 merge  place  bypass 
    -- predecessors 1619 1645 
    -- successors 1647 
    -- members (1) 
      -- 	branch_block_stmt_2042/merge_stmt_2635_PhiReqMerge
      -- 
    cp_elements(1646) <= OrReduce(cp_elements(1619) & cp_elements(1645));
    -- CP-element group 1647 fork  transition  bypass 
    -- predecessors 1646 
    -- successors 1648 1649 
    -- members (1) 
      -- 	branch_block_stmt_2042/merge_stmt_2635_PhiAck/$entry
      -- 
    cp_elements(1647) <= cp_elements(1646);
    -- CP-element group 1648 transition  input  bypass 
    -- predecessors 1647 
    -- successors 1650 
    -- members (1) 
      -- 	branch_block_stmt_2042/merge_stmt_2635_PhiAck/phi_stmt_2636_ack
      -- 
    phi_stmt_2636_ack_17073_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2636_ack_0, ack => cp_elements(1648)); -- 
    -- CP-element group 1649 transition  input  bypass 
    -- predecessors 1647 
    -- successors 1650 
    -- members (1) 
      -- 	branch_block_stmt_2042/merge_stmt_2635_PhiAck/phi_stmt_2642_ack
      -- 
    phi_stmt_2642_ack_17074_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2642_ack_0, ack => cp_elements(1649)); -- 
    -- CP-element group 1650 join  transition  bypass 
    -- predecessors 1648 1649 
    -- successors 25 
    -- members (1) 
      -- 	branch_block_stmt_2042/merge_stmt_2635_PhiAck/$exit
      -- 
    cp_element_group_1650: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1650"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1648) & cp_elements(1649);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1650), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1651 transition  bypass 
    -- predecessors 277 
    -- successors 1653 
    -- members (4) 
      -- 	branch_block_stmt_2042/bb_13_rotor_flux_calcx_xexit_PhiReq/phi_stmt_2683/phi_stmt_2683_sources/type_cast_2686/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_2042/bb_13_rotor_flux_calcx_xexit_PhiReq/phi_stmt_2683/phi_stmt_2683_sources/type_cast_2686/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_2042/bb_13_rotor_flux_calcx_xexit_PhiReq/phi_stmt_2683/phi_stmt_2683_sources/type_cast_2686/SplitProtocol/Sample/rr
      -- 	branch_block_stmt_2042/bb_13_rotor_flux_calcx_xexit_PhiReq/phi_stmt_2683/phi_stmt_2683_sources/type_cast_2686/SplitProtocol/Sample/ra
      -- 
    cp_elements(1651) <= cp_elements(277);
    -- CP-element group 1652 transition  bypass 
    -- predecessors 277 
    -- successors 1653 
    -- members (4) 
      -- 	branch_block_stmt_2042/bb_13_rotor_flux_calcx_xexit_PhiReq/phi_stmt_2683/phi_stmt_2683_sources/type_cast_2686/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_2042/bb_13_rotor_flux_calcx_xexit_PhiReq/phi_stmt_2683/phi_stmt_2683_sources/type_cast_2686/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_2042/bb_13_rotor_flux_calcx_xexit_PhiReq/phi_stmt_2683/phi_stmt_2683_sources/type_cast_2686/SplitProtocol/Update/cr
      -- 	branch_block_stmt_2042/bb_13_rotor_flux_calcx_xexit_PhiReq/phi_stmt_2683/phi_stmt_2683_sources/type_cast_2686/SplitProtocol/Update/ca
      -- 
    cp_elements(1652) <= cp_elements(277);
    -- CP-element group 1653 join  transition  output  bypass 
    -- predecessors 1651 1652 
    -- successors 1659 
    -- members (6) 
      -- 	branch_block_stmt_2042/bb_13_rotor_flux_calcx_xexit_PhiReq/$exit
      -- 	branch_block_stmt_2042/bb_13_rotor_flux_calcx_xexit_PhiReq/phi_stmt_2683/$exit
      -- 	branch_block_stmt_2042/bb_13_rotor_flux_calcx_xexit_PhiReq/phi_stmt_2683/phi_stmt_2683_sources/$exit
      -- 	branch_block_stmt_2042/bb_13_rotor_flux_calcx_xexit_PhiReq/phi_stmt_2683/phi_stmt_2683_sources/type_cast_2686/$exit
      -- 	branch_block_stmt_2042/bb_13_rotor_flux_calcx_xexit_PhiReq/phi_stmt_2683/phi_stmt_2683_sources/type_cast_2686/SplitProtocol/$exit
      -- 	branch_block_stmt_2042/bb_13_rotor_flux_calcx_xexit_PhiReq/phi_stmt_2683/phi_stmt_2683_req
      -- 
    cp_element_group_1653: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1653"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1651) & cp_elements(1652);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1653), clk => clk, reset => reset); --
    end block;
    phi_stmt_2683_req_17100_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1653), ack => phi_stmt_2683_req_1); -- 
    -- CP-element group 1654 transition  output  bypass 
    -- predecessors 459 
    -- successors 1655 
    -- members (2) 
      -- 	branch_block_stmt_2042/xx_xcritedgex_xix_xi52_rotor_flux_calcx_xexit_PhiReq/phi_stmt_2683/phi_stmt_2683_sources/type_cast_2686/SplitProtocol/Sample/rr
      -- 	branch_block_stmt_2042/xx_xcritedgex_xix_xi52_rotor_flux_calcx_xexit_PhiReq/phi_stmt_2683/phi_stmt_2683_sources/type_cast_2686/SplitProtocol/Sample/$entry
      -- 
    cp_elements(1654) <= cp_elements(459);
    rr_17119_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1654), ack => type_cast_2686_inst_req_0); -- 
    -- CP-element group 1655 transition  input  bypass 
    -- predecessors 1654 
    -- successors 1658 
    -- members (2) 
      -- 	branch_block_stmt_2042/xx_xcritedgex_xix_xi52_rotor_flux_calcx_xexit_PhiReq/phi_stmt_2683/phi_stmt_2683_sources/type_cast_2686/SplitProtocol/Sample/ra
      -- 	branch_block_stmt_2042/xx_xcritedgex_xix_xi52_rotor_flux_calcx_xexit_PhiReq/phi_stmt_2683/phi_stmt_2683_sources/type_cast_2686/SplitProtocol/Sample/$exit
      -- 
    ra_17120_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2686_inst_ack_0, ack => cp_elements(1655)); -- 
    -- CP-element group 1656 transition  output  bypass 
    -- predecessors 459 
    -- successors 1657 
    -- members (2) 
      -- 	branch_block_stmt_2042/xx_xcritedgex_xix_xi52_rotor_flux_calcx_xexit_PhiReq/phi_stmt_2683/phi_stmt_2683_sources/type_cast_2686/SplitProtocol/Update/cr
      -- 	branch_block_stmt_2042/xx_xcritedgex_xix_xi52_rotor_flux_calcx_xexit_PhiReq/phi_stmt_2683/phi_stmt_2683_sources/type_cast_2686/SplitProtocol/Update/$entry
      -- 
    cp_elements(1656) <= cp_elements(459);
    cr_17124_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1656), ack => type_cast_2686_inst_req_1); -- 
    -- CP-element group 1657 transition  input  bypass 
    -- predecessors 1656 
    -- successors 1658 
    -- members (2) 
      -- 	branch_block_stmt_2042/xx_xcritedgex_xix_xi52_rotor_flux_calcx_xexit_PhiReq/phi_stmt_2683/phi_stmt_2683_sources/type_cast_2686/SplitProtocol/Update/ca
      -- 	branch_block_stmt_2042/xx_xcritedgex_xix_xi52_rotor_flux_calcx_xexit_PhiReq/phi_stmt_2683/phi_stmt_2683_sources/type_cast_2686/SplitProtocol/Update/$exit
      -- 
    ca_17125_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2686_inst_ack_1, ack => cp_elements(1657)); -- 
    -- CP-element group 1658 join  transition  output  bypass 
    -- predecessors 1655 1657 
    -- successors 1659 
    -- members (6) 
      -- 	branch_block_stmt_2042/xx_xcritedgex_xix_xi52_rotor_flux_calcx_xexit_PhiReq/phi_stmt_2683/phi_stmt_2683_req
      -- 	branch_block_stmt_2042/xx_xcritedgex_xix_xi52_rotor_flux_calcx_xexit_PhiReq/phi_stmt_2683/phi_stmt_2683_sources/type_cast_2686/SplitProtocol/$exit
      -- 	branch_block_stmt_2042/xx_xcritedgex_xix_xi52_rotor_flux_calcx_xexit_PhiReq/$exit
      -- 	branch_block_stmt_2042/xx_xcritedgex_xix_xi52_rotor_flux_calcx_xexit_PhiReq/phi_stmt_2683/$exit
      -- 	branch_block_stmt_2042/xx_xcritedgex_xix_xi52_rotor_flux_calcx_xexit_PhiReq/phi_stmt_2683/phi_stmt_2683_sources/$exit
      -- 	branch_block_stmt_2042/xx_xcritedgex_xix_xi52_rotor_flux_calcx_xexit_PhiReq/phi_stmt_2683/phi_stmt_2683_sources/type_cast_2686/$exit
      -- 
    cp_element_group_1658: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1658"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1655) & cp_elements(1657);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1658), clk => clk, reset => reset); --
    end block;
    phi_stmt_2683_req_17126_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1658), ack => phi_stmt_2683_req_0); -- 
    -- CP-element group 1659 merge  place  bypass 
    -- predecessors 1653 1658 
    -- successors 1660 
    -- members (1) 
      -- 	branch_block_stmt_2042/merge_stmt_2682_PhiReqMerge
      -- 
    cp_elements(1659) <= OrReduce(cp_elements(1653) & cp_elements(1658));
    -- CP-element group 1660 transition  bypass 
    -- predecessors 1659 
    -- successors 1661 
    -- members (1) 
      -- 	branch_block_stmt_2042/merge_stmt_2682_PhiAck/$entry
      -- 
    cp_elements(1660) <= cp_elements(1659);
    -- CP-element group 1661 transition  place  input  bypass 
    -- predecessors 1660 
    -- successors 460 
    -- members (4) 
      -- 	branch_block_stmt_2042/merge_stmt_2682__exit__
      -- 	branch_block_stmt_2042/assign_stmt_2696_to_assign_stmt_2716__entry__
      -- 	branch_block_stmt_2042/merge_stmt_2682_PhiAck/phi_stmt_2683_ack
      -- 	branch_block_stmt_2042/merge_stmt_2682_PhiAck/$exit
      -- 
    phi_stmt_2683_ack_17131_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2683_ack_0, ack => cp_elements(1661)); -- 
    -- CP-element group 1662 fork  transition  bypass 
    -- predecessors 29 
    -- successors 1663 1675 
    -- members (1) 
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xix_xi5x_xpreheader_bbx_xnph7x_xix_xix_xi5_PhiReq/$entry
      -- 
    cp_elements(1662) <= cp_elements(29);
    -- CP-element group 1663 fork  transition  bypass 
    -- predecessors 1662 
    -- successors 1664 1668 
    -- members (2) 
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xix_xi5x_xpreheader_bbx_xnph7x_xix_xix_xi5_PhiReq/phi_stmt_2813/phi_stmt_2813_sources/$entry
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xix_xi5x_xpreheader_bbx_xnph7x_xix_xix_xi5_PhiReq/phi_stmt_2813/$entry
      -- 
    cp_elements(1663) <= cp_elements(1662);
    -- CP-element group 1664 fork  transition  bypass 
    -- predecessors 1663 
    -- successors 1665 1666 
    -- members (2) 
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xix_xi5x_xpreheader_bbx_xnph7x_xix_xix_xi5_PhiReq/phi_stmt_2813/phi_stmt_2813_sources/type_cast_2816/SplitProtocol/$entry
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xix_xi5x_xpreheader_bbx_xnph7x_xix_xix_xi5_PhiReq/phi_stmt_2813/phi_stmt_2813_sources/type_cast_2816/$entry
      -- 
    cp_elements(1664) <= cp_elements(1663);
    -- CP-element group 1665 transition  bypass 
    -- predecessors 1664 
    -- successors 1667 
    -- members (4) 
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xix_xi5x_xpreheader_bbx_xnph7x_xix_xix_xi5_PhiReq/phi_stmt_2813/phi_stmt_2813_sources/type_cast_2816/SplitProtocol/Sample/ra
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xix_xi5x_xpreheader_bbx_xnph7x_xix_xix_xi5_PhiReq/phi_stmt_2813/phi_stmt_2813_sources/type_cast_2816/SplitProtocol/Sample/rr
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xix_xi5x_xpreheader_bbx_xnph7x_xix_xix_xi5_PhiReq/phi_stmt_2813/phi_stmt_2813_sources/type_cast_2816/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xix_xi5x_xpreheader_bbx_xnph7x_xix_xix_xi5_PhiReq/phi_stmt_2813/phi_stmt_2813_sources/type_cast_2816/SplitProtocol/Sample/$entry
      -- 
    cp_elements(1665) <= cp_elements(1664);
    -- CP-element group 1666 transition  bypass 
    -- predecessors 1664 
    -- successors 1667 
    -- members (4) 
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xix_xi5x_xpreheader_bbx_xnph7x_xix_xix_xi5_PhiReq/phi_stmt_2813/phi_stmt_2813_sources/type_cast_2816/SplitProtocol/Update/ca
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xix_xi5x_xpreheader_bbx_xnph7x_xix_xix_xi5_PhiReq/phi_stmt_2813/phi_stmt_2813_sources/type_cast_2816/SplitProtocol/Update/cr
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xix_xi5x_xpreheader_bbx_xnph7x_xix_xix_xi5_PhiReq/phi_stmt_2813/phi_stmt_2813_sources/type_cast_2816/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xix_xi5x_xpreheader_bbx_xnph7x_xix_xix_xi5_PhiReq/phi_stmt_2813/phi_stmt_2813_sources/type_cast_2816/SplitProtocol/Update/$entry
      -- 
    cp_elements(1666) <= cp_elements(1664);
    -- CP-element group 1667 join  transition  bypass 
    -- predecessors 1665 1666 
    -- successors 1674 
    -- members (2) 
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xix_xi5x_xpreheader_bbx_xnph7x_xix_xix_xi5_PhiReq/phi_stmt_2813/phi_stmt_2813_sources/type_cast_2816/SplitProtocol/$exit
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xix_xi5x_xpreheader_bbx_xnph7x_xix_xix_xi5_PhiReq/phi_stmt_2813/phi_stmt_2813_sources/type_cast_2816/$exit
      -- 
    cp_element_group_1667: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1667"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1665) & cp_elements(1666);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1667), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1668 fork  transition  bypass 
    -- predecessors 1663 
    -- successors 1669 1671 
    -- members (2) 
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xix_xi5x_xpreheader_bbx_xnph7x_xix_xix_xi5_PhiReq/phi_stmt_2813/phi_stmt_2813_sources/type_cast_2818/SplitProtocol/$entry
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xix_xi5x_xpreheader_bbx_xnph7x_xix_xix_xi5_PhiReq/phi_stmt_2813/phi_stmt_2813_sources/type_cast_2818/$entry
      -- 
    cp_elements(1668) <= cp_elements(1663);
    -- CP-element group 1669 transition  output  bypass 
    -- predecessors 1668 
    -- successors 1670 
    -- members (2) 
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xix_xi5x_xpreheader_bbx_xnph7x_xix_xix_xi5_PhiReq/phi_stmt_2813/phi_stmt_2813_sources/type_cast_2818/SplitProtocol/Sample/rr
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xix_xi5x_xpreheader_bbx_xnph7x_xix_xix_xi5_PhiReq/phi_stmt_2813/phi_stmt_2813_sources/type_cast_2818/SplitProtocol/Sample/$entry
      -- 
    cp_elements(1669) <= cp_elements(1668);
    rr_17190_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1669), ack => type_cast_2818_inst_req_0); -- 
    -- CP-element group 1670 transition  input  bypass 
    -- predecessors 1669 
    -- successors 1673 
    -- members (2) 
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xix_xi5x_xpreheader_bbx_xnph7x_xix_xix_xi5_PhiReq/phi_stmt_2813/phi_stmt_2813_sources/type_cast_2818/SplitProtocol/Sample/ra
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xix_xi5x_xpreheader_bbx_xnph7x_xix_xix_xi5_PhiReq/phi_stmt_2813/phi_stmt_2813_sources/type_cast_2818/SplitProtocol/Sample/$exit
      -- 
    ra_17191_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2818_inst_ack_0, ack => cp_elements(1670)); -- 
    -- CP-element group 1671 transition  output  bypass 
    -- predecessors 1668 
    -- successors 1672 
    -- members (2) 
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xix_xi5x_xpreheader_bbx_xnph7x_xix_xix_xi5_PhiReq/phi_stmt_2813/phi_stmt_2813_sources/type_cast_2818/SplitProtocol/Update/cr
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xix_xi5x_xpreheader_bbx_xnph7x_xix_xix_xi5_PhiReq/phi_stmt_2813/phi_stmt_2813_sources/type_cast_2818/SplitProtocol/Update/$entry
      -- 
    cp_elements(1671) <= cp_elements(1668);
    cr_17195_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1671), ack => type_cast_2818_inst_req_1); -- 
    -- CP-element group 1672 transition  input  bypass 
    -- predecessors 1671 
    -- successors 1673 
    -- members (2) 
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xix_xi5x_xpreheader_bbx_xnph7x_xix_xix_xi5_PhiReq/phi_stmt_2813/phi_stmt_2813_sources/type_cast_2818/SplitProtocol/Update/ca
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xix_xi5x_xpreheader_bbx_xnph7x_xix_xix_xi5_PhiReq/phi_stmt_2813/phi_stmt_2813_sources/type_cast_2818/SplitProtocol/Update/$exit
      -- 
    ca_17196_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2818_inst_ack_1, ack => cp_elements(1672)); -- 
    -- CP-element group 1673 join  transition  bypass 
    -- predecessors 1670 1672 
    -- successors 1674 
    -- members (2) 
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xix_xi5x_xpreheader_bbx_xnph7x_xix_xix_xi5_PhiReq/phi_stmt_2813/phi_stmt_2813_sources/type_cast_2818/SplitProtocol/$exit
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xix_xi5x_xpreheader_bbx_xnph7x_xix_xix_xi5_PhiReq/phi_stmt_2813/phi_stmt_2813_sources/type_cast_2818/$exit
      -- 
    cp_element_group_1673: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1673"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1670) & cp_elements(1672);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1673), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1674 join  transition  output  bypass 
    -- predecessors 1667 1673 
    -- successors 1679 
    -- members (3) 
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xix_xi5x_xpreheader_bbx_xnph7x_xix_xix_xi5_PhiReq/phi_stmt_2813/phi_stmt_2813_req
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xix_xi5x_xpreheader_bbx_xnph7x_xix_xix_xi5_PhiReq/phi_stmt_2813/phi_stmt_2813_sources/$exit
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xix_xi5x_xpreheader_bbx_xnph7x_xix_xix_xi5_PhiReq/phi_stmt_2813/$exit
      -- 
    cp_element_group_1674: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1674"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1667) & cp_elements(1673);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1674), clk => clk, reset => reset); --
    end block;
    phi_stmt_2813_req_17197_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1674), ack => phi_stmt_2813_req_1); -- 
    -- CP-element group 1675 fork  transition  bypass 
    -- predecessors 1662 
    -- successors 1676 1677 
    -- members (4) 
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xix_xi5x_xpreheader_bbx_xnph7x_xix_xix_xi5_PhiReq/phi_stmt_2819/phi_stmt_2819_sources/type_cast_2822/SplitProtocol/$entry
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xix_xi5x_xpreheader_bbx_xnph7x_xix_xix_xi5_PhiReq/phi_stmt_2819/phi_stmt_2819_sources/type_cast_2822/$entry
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xix_xi5x_xpreheader_bbx_xnph7x_xix_xix_xi5_PhiReq/phi_stmt_2819/phi_stmt_2819_sources/$entry
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xix_xi5x_xpreheader_bbx_xnph7x_xix_xix_xi5_PhiReq/phi_stmt_2819/$entry
      -- 
    cp_elements(1675) <= cp_elements(1662);
    -- CP-element group 1676 transition  bypass 
    -- predecessors 1675 
    -- successors 1678 
    -- members (4) 
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xix_xi5x_xpreheader_bbx_xnph7x_xix_xix_xi5_PhiReq/phi_stmt_2819/phi_stmt_2819_sources/type_cast_2822/SplitProtocol/Sample/ra
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xix_xi5x_xpreheader_bbx_xnph7x_xix_xix_xi5_PhiReq/phi_stmt_2819/phi_stmt_2819_sources/type_cast_2822/SplitProtocol/Sample/rr
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xix_xi5x_xpreheader_bbx_xnph7x_xix_xix_xi5_PhiReq/phi_stmt_2819/phi_stmt_2819_sources/type_cast_2822/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xix_xi5x_xpreheader_bbx_xnph7x_xix_xix_xi5_PhiReq/phi_stmt_2819/phi_stmt_2819_sources/type_cast_2822/SplitProtocol/Sample/$entry
      -- 
    cp_elements(1676) <= cp_elements(1675);
    -- CP-element group 1677 transition  bypass 
    -- predecessors 1675 
    -- successors 1678 
    -- members (4) 
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xix_xi5x_xpreheader_bbx_xnph7x_xix_xix_xi5_PhiReq/phi_stmt_2819/phi_stmt_2819_sources/type_cast_2822/SplitProtocol/Update/ca
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xix_xi5x_xpreheader_bbx_xnph7x_xix_xix_xi5_PhiReq/phi_stmt_2819/phi_stmt_2819_sources/type_cast_2822/SplitProtocol/Update/cr
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xix_xi5x_xpreheader_bbx_xnph7x_xix_xix_xi5_PhiReq/phi_stmt_2819/phi_stmt_2819_sources/type_cast_2822/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xix_xi5x_xpreheader_bbx_xnph7x_xix_xix_xi5_PhiReq/phi_stmt_2819/phi_stmt_2819_sources/type_cast_2822/SplitProtocol/Update/$entry
      -- 
    cp_elements(1677) <= cp_elements(1675);
    -- CP-element group 1678 join  transition  output  bypass 
    -- predecessors 1676 1677 
    -- successors 1679 
    -- members (5) 
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xix_xi5x_xpreheader_bbx_xnph7x_xix_xix_xi5_PhiReq/phi_stmt_2819/phi_stmt_2819_req
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xix_xi5x_xpreheader_bbx_xnph7x_xix_xix_xi5_PhiReq/phi_stmt_2819/phi_stmt_2819_sources/type_cast_2822/SplitProtocol/$exit
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xix_xi5x_xpreheader_bbx_xnph7x_xix_xix_xi5_PhiReq/phi_stmt_2819/phi_stmt_2819_sources/type_cast_2822/$exit
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xix_xi5x_xpreheader_bbx_xnph7x_xix_xix_xi5_PhiReq/phi_stmt_2819/phi_stmt_2819_sources/$exit
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xix_xi5x_xpreheader_bbx_xnph7x_xix_xix_xi5_PhiReq/phi_stmt_2819/$exit
      -- 
    cp_element_group_1678: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1678"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1676) & cp_elements(1677);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1678), clk => clk, reset => reset); --
    end block;
    phi_stmt_2819_req_17220_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1678), ack => phi_stmt_2819_req_1); -- 
    -- CP-element group 1679 join  transition  bypass 
    -- predecessors 1674 1678 
    -- successors 1700 
    -- members (1) 
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xix_xi5x_xpreheader_bbx_xnph7x_xix_xix_xi5_PhiReq/$exit
      -- 
    cp_element_group_1679: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1679"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1674) & cp_elements(1678);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1679), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1680 fork  transition  bypass 
    -- predecessors 624 
    -- successors 1681 1693 
    -- members (1) 
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi11_bbx_xnph7x_xix_xix_xi5_PhiReq/$entry
      -- 
    cp_elements(1680) <= cp_elements(624);
    -- CP-element group 1681 fork  transition  bypass 
    -- predecessors 1680 
    -- successors 1682 1688 
    -- members (2) 
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi11_bbx_xnph7x_xix_xix_xi5_PhiReq/phi_stmt_2813/phi_stmt_2813_sources/$entry
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi11_bbx_xnph7x_xix_xix_xi5_PhiReq/phi_stmt_2813/$entry
      -- 
    cp_elements(1681) <= cp_elements(1680);
    -- CP-element group 1682 fork  transition  bypass 
    -- predecessors 1681 
    -- successors 1683 1685 
    -- members (2) 
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi11_bbx_xnph7x_xix_xix_xi5_PhiReq/phi_stmt_2813/phi_stmt_2813_sources/type_cast_2816/SplitProtocol/$entry
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi11_bbx_xnph7x_xix_xix_xi5_PhiReq/phi_stmt_2813/phi_stmt_2813_sources/type_cast_2816/$entry
      -- 
    cp_elements(1682) <= cp_elements(1681);
    -- CP-element group 1683 transition  output  bypass 
    -- predecessors 1682 
    -- successors 1684 
    -- members (2) 
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi11_bbx_xnph7x_xix_xix_xi5_PhiReq/phi_stmt_2813/phi_stmt_2813_sources/type_cast_2816/SplitProtocol/Sample/rr
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi11_bbx_xnph7x_xix_xix_xi5_PhiReq/phi_stmt_2813/phi_stmt_2813_sources/type_cast_2816/SplitProtocol/Sample/$entry
      -- 
    cp_elements(1683) <= cp_elements(1682);
    rr_17239_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1683), ack => type_cast_2816_inst_req_0); -- 
    -- CP-element group 1684 transition  input  bypass 
    -- predecessors 1683 
    -- successors 1687 
    -- members (2) 
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi11_bbx_xnph7x_xix_xix_xi5_PhiReq/phi_stmt_2813/phi_stmt_2813_sources/type_cast_2816/SplitProtocol/Sample/ra
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi11_bbx_xnph7x_xix_xix_xi5_PhiReq/phi_stmt_2813/phi_stmt_2813_sources/type_cast_2816/SplitProtocol/Sample/$exit
      -- 
    ra_17240_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2816_inst_ack_0, ack => cp_elements(1684)); -- 
    -- CP-element group 1685 transition  output  bypass 
    -- predecessors 1682 
    -- successors 1686 
    -- members (2) 
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi11_bbx_xnph7x_xix_xix_xi5_PhiReq/phi_stmt_2813/phi_stmt_2813_sources/type_cast_2816/SplitProtocol/Update/cr
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi11_bbx_xnph7x_xix_xix_xi5_PhiReq/phi_stmt_2813/phi_stmt_2813_sources/type_cast_2816/SplitProtocol/Update/$entry
      -- 
    cp_elements(1685) <= cp_elements(1682);
    cr_17244_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1685), ack => type_cast_2816_inst_req_1); -- 
    -- CP-element group 1686 transition  input  bypass 
    -- predecessors 1685 
    -- successors 1687 
    -- members (2) 
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi11_bbx_xnph7x_xix_xix_xi5_PhiReq/phi_stmt_2813/phi_stmt_2813_sources/type_cast_2816/SplitProtocol/Update/ca
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi11_bbx_xnph7x_xix_xix_xi5_PhiReq/phi_stmt_2813/phi_stmt_2813_sources/type_cast_2816/SplitProtocol/Update/$exit
      -- 
    ca_17245_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2816_inst_ack_1, ack => cp_elements(1686)); -- 
    -- CP-element group 1687 join  transition  bypass 
    -- predecessors 1684 1686 
    -- successors 1692 
    -- members (2) 
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi11_bbx_xnph7x_xix_xix_xi5_PhiReq/phi_stmt_2813/phi_stmt_2813_sources/type_cast_2816/SplitProtocol/$exit
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi11_bbx_xnph7x_xix_xix_xi5_PhiReq/phi_stmt_2813/phi_stmt_2813_sources/type_cast_2816/$exit
      -- 
    cp_element_group_1687: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1687"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1684) & cp_elements(1686);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1687), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1688 fork  transition  bypass 
    -- predecessors 1681 
    -- successors 1689 1690 
    -- members (2) 
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi11_bbx_xnph7x_xix_xix_xi5_PhiReq/phi_stmt_2813/phi_stmt_2813_sources/type_cast_2818/$entry
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi11_bbx_xnph7x_xix_xix_xi5_PhiReq/phi_stmt_2813/phi_stmt_2813_sources/type_cast_2818/SplitProtocol/$entry
      -- 
    cp_elements(1688) <= cp_elements(1681);
    -- CP-element group 1689 transition  bypass 
    -- predecessors 1688 
    -- successors 1691 
    -- members (4) 
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi11_bbx_xnph7x_xix_xix_xi5_PhiReq/phi_stmt_2813/phi_stmt_2813_sources/type_cast_2818/SplitProtocol/Sample/ra
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi11_bbx_xnph7x_xix_xix_xi5_PhiReq/phi_stmt_2813/phi_stmt_2813_sources/type_cast_2818/SplitProtocol/Sample/rr
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi11_bbx_xnph7x_xix_xix_xi5_PhiReq/phi_stmt_2813/phi_stmt_2813_sources/type_cast_2818/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi11_bbx_xnph7x_xix_xix_xi5_PhiReq/phi_stmt_2813/phi_stmt_2813_sources/type_cast_2818/SplitProtocol/Sample/$entry
      -- 
    cp_elements(1689) <= cp_elements(1688);
    -- CP-element group 1690 transition  bypass 
    -- predecessors 1688 
    -- successors 1691 
    -- members (4) 
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi11_bbx_xnph7x_xix_xix_xi5_PhiReq/phi_stmt_2813/phi_stmt_2813_sources/type_cast_2818/SplitProtocol/Update/ca
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi11_bbx_xnph7x_xix_xix_xi5_PhiReq/phi_stmt_2813/phi_stmt_2813_sources/type_cast_2818/SplitProtocol/Update/cr
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi11_bbx_xnph7x_xix_xix_xi5_PhiReq/phi_stmt_2813/phi_stmt_2813_sources/type_cast_2818/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi11_bbx_xnph7x_xix_xix_xi5_PhiReq/phi_stmt_2813/phi_stmt_2813_sources/type_cast_2818/SplitProtocol/Update/$entry
      -- 
    cp_elements(1690) <= cp_elements(1688);
    -- CP-element group 1691 join  transition  bypass 
    -- predecessors 1689 1690 
    -- successors 1692 
    -- members (2) 
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi11_bbx_xnph7x_xix_xix_xi5_PhiReq/phi_stmt_2813/phi_stmt_2813_sources/type_cast_2818/SplitProtocol/$exit
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi11_bbx_xnph7x_xix_xix_xi5_PhiReq/phi_stmt_2813/phi_stmt_2813_sources/type_cast_2818/$exit
      -- 
    cp_element_group_1691: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1691"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1689) & cp_elements(1690);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1691), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1692 join  transition  output  bypass 
    -- predecessors 1687 1691 
    -- successors 1699 
    -- members (3) 
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi11_bbx_xnph7x_xix_xix_xi5_PhiReq/phi_stmt_2813/phi_stmt_2813_req
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi11_bbx_xnph7x_xix_xix_xi5_PhiReq/phi_stmt_2813/phi_stmt_2813_sources/$exit
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi11_bbx_xnph7x_xix_xix_xi5_PhiReq/phi_stmt_2813/$exit
      -- 
    cp_element_group_1692: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1692"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1687) & cp_elements(1691);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1692), clk => clk, reset => reset); --
    end block;
    phi_stmt_2813_req_17262_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1692), ack => phi_stmt_2813_req_0); -- 
    -- CP-element group 1693 fork  transition  bypass 
    -- predecessors 1680 
    -- successors 1694 1696 
    -- members (4) 
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi11_bbx_xnph7x_xix_xix_xi5_PhiReq/phi_stmt_2819/$entry
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi11_bbx_xnph7x_xix_xix_xi5_PhiReq/phi_stmt_2819/phi_stmt_2819_sources/$entry
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi11_bbx_xnph7x_xix_xix_xi5_PhiReq/phi_stmt_2819/phi_stmt_2819_sources/type_cast_2822/$entry
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi11_bbx_xnph7x_xix_xix_xi5_PhiReq/phi_stmt_2819/phi_stmt_2819_sources/type_cast_2822/SplitProtocol/$entry
      -- 
    cp_elements(1693) <= cp_elements(1680);
    -- CP-element group 1694 transition  output  bypass 
    -- predecessors 1693 
    -- successors 1695 
    -- members (2) 
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi11_bbx_xnph7x_xix_xix_xi5_PhiReq/phi_stmt_2819/phi_stmt_2819_sources/type_cast_2822/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi11_bbx_xnph7x_xix_xix_xi5_PhiReq/phi_stmt_2819/phi_stmt_2819_sources/type_cast_2822/SplitProtocol/Sample/rr
      -- 
    cp_elements(1694) <= cp_elements(1693);
    rr_17278_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1694), ack => type_cast_2822_inst_req_0); -- 
    -- CP-element group 1695 transition  input  bypass 
    -- predecessors 1694 
    -- successors 1698 
    -- members (2) 
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi11_bbx_xnph7x_xix_xix_xi5_PhiReq/phi_stmt_2819/phi_stmt_2819_sources/type_cast_2822/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi11_bbx_xnph7x_xix_xix_xi5_PhiReq/phi_stmt_2819/phi_stmt_2819_sources/type_cast_2822/SplitProtocol/Sample/ra
      -- 
    ra_17279_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2822_inst_ack_0, ack => cp_elements(1695)); -- 
    -- CP-element group 1696 transition  output  bypass 
    -- predecessors 1693 
    -- successors 1697 
    -- members (2) 
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi11_bbx_xnph7x_xix_xix_xi5_PhiReq/phi_stmt_2819/phi_stmt_2819_sources/type_cast_2822/SplitProtocol/Update/cr
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi11_bbx_xnph7x_xix_xix_xi5_PhiReq/phi_stmt_2819/phi_stmt_2819_sources/type_cast_2822/SplitProtocol/Update/$entry
      -- 
    cp_elements(1696) <= cp_elements(1693);
    cr_17283_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1696), ack => type_cast_2822_inst_req_1); -- 
    -- CP-element group 1697 transition  input  bypass 
    -- predecessors 1696 
    -- successors 1698 
    -- members (2) 
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi11_bbx_xnph7x_xix_xix_xi5_PhiReq/phi_stmt_2819/phi_stmt_2819_sources/type_cast_2822/SplitProtocol/Update/ca
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi11_bbx_xnph7x_xix_xix_xi5_PhiReq/phi_stmt_2819/phi_stmt_2819_sources/type_cast_2822/SplitProtocol/Update/$exit
      -- 
    ca_17284_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2822_inst_ack_1, ack => cp_elements(1697)); -- 
    -- CP-element group 1698 join  transition  output  bypass 
    -- predecessors 1695 1697 
    -- successors 1699 
    -- members (5) 
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi11_bbx_xnph7x_xix_xix_xi5_PhiReq/phi_stmt_2819/phi_stmt_2819_req
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi11_bbx_xnph7x_xix_xix_xi5_PhiReq/phi_stmt_2819/phi_stmt_2819_sources/type_cast_2822/SplitProtocol/$exit
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi11_bbx_xnph7x_xix_xix_xi5_PhiReq/phi_stmt_2819/phi_stmt_2819_sources/type_cast_2822/$exit
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi11_bbx_xnph7x_xix_xix_xi5_PhiReq/phi_stmt_2819/phi_stmt_2819_sources/$exit
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi11_bbx_xnph7x_xix_xix_xi5_PhiReq/phi_stmt_2819/$exit
      -- 
    cp_element_group_1698: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1698"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1695) & cp_elements(1697);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1698), clk => clk, reset => reset); --
    end block;
    phi_stmt_2819_req_17285_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1698), ack => phi_stmt_2819_req_0); -- 
    -- CP-element group 1699 join  transition  bypass 
    -- predecessors 1692 1698 
    -- successors 1700 
    -- members (1) 
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi11_bbx_xnph7x_xix_xix_xi5_PhiReq/$exit
      -- 
    cp_element_group_1699: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1699"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1692) & cp_elements(1698);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1699), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1700 merge  place  bypass 
    -- predecessors 1679 1699 
    -- successors 1701 
    -- members (1) 
      -- 	branch_block_stmt_2042/merge_stmt_2812_PhiReqMerge
      -- 
    cp_elements(1700) <= OrReduce(cp_elements(1679) & cp_elements(1699));
    -- CP-element group 1701 fork  transition  bypass 
    -- predecessors 1700 
    -- successors 1702 1703 
    -- members (1) 
      -- 	branch_block_stmt_2042/merge_stmt_2812_PhiAck/$entry
      -- 
    cp_elements(1701) <= cp_elements(1700);
    -- CP-element group 1702 transition  input  bypass 
    -- predecessors 1701 
    -- successors 1704 
    -- members (1) 
      -- 	branch_block_stmt_2042/merge_stmt_2812_PhiAck/phi_stmt_2813_ack
      -- 
    phi_stmt_2813_ack_17290_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2813_ack_0, ack => cp_elements(1702)); -- 
    -- CP-element group 1703 transition  input  bypass 
    -- predecessors 1701 
    -- successors 1704 
    -- members (1) 
      -- 	branch_block_stmt_2042/merge_stmt_2812_PhiAck/phi_stmt_2819_ack
      -- 
    phi_stmt_2819_ack_17291_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2819_ack_0, ack => cp_elements(1703)); -- 
    -- CP-element group 1704 join  transition  bypass 
    -- predecessors 1702 1703 
    -- successors 30 
    -- members (1) 
      -- 	branch_block_stmt_2042/merge_stmt_2812_PhiAck/$exit
      -- 
    cp_element_group_1704: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1704"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1702) & cp_elements(1703);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1704), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1705 fork  transition  bypass 
    -- predecessors 596 
    -- successors 1706 1718 
    -- members (1) 
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi8_bbx_xnphx_xix_xix_xi8_PhiReq/$entry
      -- 
    cp_elements(1705) <= cp_elements(596);
    -- CP-element group 1706 fork  transition  bypass 
    -- predecessors 1705 
    -- successors 1707 1713 
    -- members (2) 
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi8_bbx_xnphx_xix_xix_xi8_PhiReq/phi_stmt_2847/$entry
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi8_bbx_xnphx_xix_xix_xi8_PhiReq/phi_stmt_2847/phi_stmt_2847_sources/$entry
      -- 
    cp_elements(1706) <= cp_elements(1705);
    -- CP-element group 1707 fork  transition  bypass 
    -- predecessors 1706 
    -- successors 1708 1710 
    -- members (2) 
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi8_bbx_xnphx_xix_xix_xi8_PhiReq/phi_stmt_2847/phi_stmt_2847_sources/type_cast_2850/$entry
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi8_bbx_xnphx_xix_xix_xi8_PhiReq/phi_stmt_2847/phi_stmt_2847_sources/type_cast_2850/SplitProtocol/$entry
      -- 
    cp_elements(1707) <= cp_elements(1706);
    -- CP-element group 1708 transition  output  bypass 
    -- predecessors 1707 
    -- successors 1709 
    -- members (2) 
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi8_bbx_xnphx_xix_xix_xi8_PhiReq/phi_stmt_2847/phi_stmt_2847_sources/type_cast_2850/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi8_bbx_xnphx_xix_xix_xi8_PhiReq/phi_stmt_2847/phi_stmt_2847_sources/type_cast_2850/SplitProtocol/Sample/rr
      -- 
    cp_elements(1708) <= cp_elements(1707);
    rr_17322_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1708), ack => type_cast_2850_inst_req_0); -- 
    -- CP-element group 1709 transition  input  bypass 
    -- predecessors 1708 
    -- successors 1712 
    -- members (2) 
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi8_bbx_xnphx_xix_xix_xi8_PhiReq/phi_stmt_2847/phi_stmt_2847_sources/type_cast_2850/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi8_bbx_xnphx_xix_xix_xi8_PhiReq/phi_stmt_2847/phi_stmt_2847_sources/type_cast_2850/SplitProtocol/Sample/ra
      -- 
    ra_17323_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2850_inst_ack_0, ack => cp_elements(1709)); -- 
    -- CP-element group 1710 transition  output  bypass 
    -- predecessors 1707 
    -- successors 1711 
    -- members (2) 
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi8_bbx_xnphx_xix_xix_xi8_PhiReq/phi_stmt_2847/phi_stmt_2847_sources/type_cast_2850/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi8_bbx_xnphx_xix_xix_xi8_PhiReq/phi_stmt_2847/phi_stmt_2847_sources/type_cast_2850/SplitProtocol/Update/cr
      -- 
    cp_elements(1710) <= cp_elements(1707);
    cr_17327_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1710), ack => type_cast_2850_inst_req_1); -- 
    -- CP-element group 1711 transition  input  bypass 
    -- predecessors 1710 
    -- successors 1712 
    -- members (2) 
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi8_bbx_xnphx_xix_xix_xi8_PhiReq/phi_stmt_2847/phi_stmt_2847_sources/type_cast_2850/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi8_bbx_xnphx_xix_xix_xi8_PhiReq/phi_stmt_2847/phi_stmt_2847_sources/type_cast_2850/SplitProtocol/Update/ca
      -- 
    ca_17328_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2850_inst_ack_1, ack => cp_elements(1711)); -- 
    -- CP-element group 1712 join  transition  bypass 
    -- predecessors 1709 1711 
    -- successors 1717 
    -- members (2) 
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi8_bbx_xnphx_xix_xix_xi8_PhiReq/phi_stmt_2847/phi_stmt_2847_sources/type_cast_2850/$exit
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi8_bbx_xnphx_xix_xix_xi8_PhiReq/phi_stmt_2847/phi_stmt_2847_sources/type_cast_2850/SplitProtocol/$exit
      -- 
    cp_element_group_1712: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1712"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1709) & cp_elements(1711);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1712), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1713 fork  transition  bypass 
    -- predecessors 1706 
    -- successors 1714 1715 
    -- members (2) 
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi8_bbx_xnphx_xix_xix_xi8_PhiReq/phi_stmt_2847/phi_stmt_2847_sources/type_cast_2852/$entry
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi8_bbx_xnphx_xix_xix_xi8_PhiReq/phi_stmt_2847/phi_stmt_2847_sources/type_cast_2852/SplitProtocol/$entry
      -- 
    cp_elements(1713) <= cp_elements(1706);
    -- CP-element group 1714 transition  bypass 
    -- predecessors 1713 
    -- successors 1716 
    -- members (4) 
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi8_bbx_xnphx_xix_xix_xi8_PhiReq/phi_stmt_2847/phi_stmt_2847_sources/type_cast_2852/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi8_bbx_xnphx_xix_xix_xi8_PhiReq/phi_stmt_2847/phi_stmt_2847_sources/type_cast_2852/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi8_bbx_xnphx_xix_xix_xi8_PhiReq/phi_stmt_2847/phi_stmt_2847_sources/type_cast_2852/SplitProtocol/Sample/rr
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi8_bbx_xnphx_xix_xix_xi8_PhiReq/phi_stmt_2847/phi_stmt_2847_sources/type_cast_2852/SplitProtocol/Sample/ra
      -- 
    cp_elements(1714) <= cp_elements(1713);
    -- CP-element group 1715 transition  bypass 
    -- predecessors 1713 
    -- successors 1716 
    -- members (4) 
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi8_bbx_xnphx_xix_xix_xi8_PhiReq/phi_stmt_2847/phi_stmt_2847_sources/type_cast_2852/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi8_bbx_xnphx_xix_xix_xi8_PhiReq/phi_stmt_2847/phi_stmt_2847_sources/type_cast_2852/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi8_bbx_xnphx_xix_xix_xi8_PhiReq/phi_stmt_2847/phi_stmt_2847_sources/type_cast_2852/SplitProtocol/Update/cr
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi8_bbx_xnphx_xix_xix_xi8_PhiReq/phi_stmt_2847/phi_stmt_2847_sources/type_cast_2852/SplitProtocol/Update/ca
      -- 
    cp_elements(1715) <= cp_elements(1713);
    -- CP-element group 1716 join  transition  bypass 
    -- predecessors 1714 1715 
    -- successors 1717 
    -- members (2) 
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi8_bbx_xnphx_xix_xix_xi8_PhiReq/phi_stmt_2847/phi_stmt_2847_sources/type_cast_2852/$exit
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi8_bbx_xnphx_xix_xix_xi8_PhiReq/phi_stmt_2847/phi_stmt_2847_sources/type_cast_2852/SplitProtocol/$exit
      -- 
    cp_element_group_1716: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1716"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1714) & cp_elements(1715);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1716), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1717 join  transition  output  bypass 
    -- predecessors 1712 1716 
    -- successors 1724 
    -- members (3) 
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi8_bbx_xnphx_xix_xix_xi8_PhiReq/phi_stmt_2847/$exit
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi8_bbx_xnphx_xix_xix_xi8_PhiReq/phi_stmt_2847/phi_stmt_2847_sources/$exit
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi8_bbx_xnphx_xix_xix_xi8_PhiReq/phi_stmt_2847/phi_stmt_2847_req
      -- 
    cp_element_group_1717: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1717"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1712) & cp_elements(1716);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1717), clk => clk, reset => reset); --
    end block;
    phi_stmt_2847_req_17345_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1717), ack => phi_stmt_2847_req_0); -- 
    -- CP-element group 1718 fork  transition  bypass 
    -- predecessors 1705 
    -- successors 1719 1721 
    -- members (4) 
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi8_bbx_xnphx_xix_xix_xi8_PhiReq/phi_stmt_2853/$entry
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi8_bbx_xnphx_xix_xix_xi8_PhiReq/phi_stmt_2853/phi_stmt_2853_sources/$entry
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi8_bbx_xnphx_xix_xix_xi8_PhiReq/phi_stmt_2853/phi_stmt_2853_sources/type_cast_2856/$entry
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi8_bbx_xnphx_xix_xix_xi8_PhiReq/phi_stmt_2853/phi_stmt_2853_sources/type_cast_2856/SplitProtocol/$entry
      -- 
    cp_elements(1718) <= cp_elements(1705);
    -- CP-element group 1719 transition  output  bypass 
    -- predecessors 1718 
    -- successors 1720 
    -- members (2) 
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi8_bbx_xnphx_xix_xix_xi8_PhiReq/phi_stmt_2853/phi_stmt_2853_sources/type_cast_2856/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi8_bbx_xnphx_xix_xix_xi8_PhiReq/phi_stmt_2853/phi_stmt_2853_sources/type_cast_2856/SplitProtocol/Sample/rr
      -- 
    cp_elements(1719) <= cp_elements(1718);
    rr_17361_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1719), ack => type_cast_2856_inst_req_0); -- 
    -- CP-element group 1720 transition  input  bypass 
    -- predecessors 1719 
    -- successors 1723 
    -- members (2) 
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi8_bbx_xnphx_xix_xix_xi8_PhiReq/phi_stmt_2853/phi_stmt_2853_sources/type_cast_2856/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi8_bbx_xnphx_xix_xix_xi8_PhiReq/phi_stmt_2853/phi_stmt_2853_sources/type_cast_2856/SplitProtocol/Sample/ra
      -- 
    ra_17362_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2856_inst_ack_0, ack => cp_elements(1720)); -- 
    -- CP-element group 1721 transition  output  bypass 
    -- predecessors 1718 
    -- successors 1722 
    -- members (2) 
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi8_bbx_xnphx_xix_xix_xi8_PhiReq/phi_stmt_2853/phi_stmt_2853_sources/type_cast_2856/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi8_bbx_xnphx_xix_xix_xi8_PhiReq/phi_stmt_2853/phi_stmt_2853_sources/type_cast_2856/SplitProtocol/Update/cr
      -- 
    cp_elements(1721) <= cp_elements(1718);
    cr_17366_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1721), ack => type_cast_2856_inst_req_1); -- 
    -- CP-element group 1722 transition  input  bypass 
    -- predecessors 1721 
    -- successors 1723 
    -- members (2) 
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi8_bbx_xnphx_xix_xix_xi8_PhiReq/phi_stmt_2853/phi_stmt_2853_sources/type_cast_2856/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi8_bbx_xnphx_xix_xix_xi8_PhiReq/phi_stmt_2853/phi_stmt_2853_sources/type_cast_2856/SplitProtocol/Update/ca
      -- 
    ca_17367_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2856_inst_ack_1, ack => cp_elements(1722)); -- 
    -- CP-element group 1723 join  transition  output  bypass 
    -- predecessors 1720 1722 
    -- successors 1724 
    -- members (5) 
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi8_bbx_xnphx_xix_xix_xi8_PhiReq/phi_stmt_2853/$exit
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi8_bbx_xnphx_xix_xix_xi8_PhiReq/phi_stmt_2853/phi_stmt_2853_sources/$exit
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi8_bbx_xnphx_xix_xix_xi8_PhiReq/phi_stmt_2853/phi_stmt_2853_sources/type_cast_2856/$exit
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi8_bbx_xnphx_xix_xix_xi8_PhiReq/phi_stmt_2853/phi_stmt_2853_sources/type_cast_2856/SplitProtocol/$exit
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi8_bbx_xnphx_xix_xix_xi8_PhiReq/phi_stmt_2853/phi_stmt_2853_req
      -- 
    cp_element_group_1723: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1723"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1720) & cp_elements(1722);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1723), clk => clk, reset => reset); --
    end block;
    phi_stmt_2853_req_17368_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1723), ack => phi_stmt_2853_req_0); -- 
    -- CP-element group 1724 join  transition  bypass 
    -- predecessors 1717 1723 
    -- successors 1743 
    -- members (1) 
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi8_bbx_xnphx_xix_xix_xi8_PhiReq/$exit
      -- 
    cp_element_group_1724: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1724"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1717) & cp_elements(1723);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1724), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1725 fork  transition  bypass 
    -- predecessors 31 
    -- successors 1726 1738 
    -- members (1) 
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi8x_xpreheader_bbx_xnphx_xix_xix_xi8_PhiReq/$entry
      -- 
    cp_elements(1725) <= cp_elements(31);
    -- CP-element group 1726 fork  transition  bypass 
    -- predecessors 1725 
    -- successors 1727 1731 
    -- members (2) 
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi8x_xpreheader_bbx_xnphx_xix_xix_xi8_PhiReq/phi_stmt_2847/$entry
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi8x_xpreheader_bbx_xnphx_xix_xix_xi8_PhiReq/phi_stmt_2847/phi_stmt_2847_sources/$entry
      -- 
    cp_elements(1726) <= cp_elements(1725);
    -- CP-element group 1727 fork  transition  bypass 
    -- predecessors 1726 
    -- successors 1728 1729 
    -- members (2) 
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi8x_xpreheader_bbx_xnphx_xix_xix_xi8_PhiReq/phi_stmt_2847/phi_stmt_2847_sources/type_cast_2850/$entry
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi8x_xpreheader_bbx_xnphx_xix_xix_xi8_PhiReq/phi_stmt_2847/phi_stmt_2847_sources/type_cast_2850/SplitProtocol/$entry
      -- 
    cp_elements(1727) <= cp_elements(1726);
    -- CP-element group 1728 transition  bypass 
    -- predecessors 1727 
    -- successors 1730 
    -- members (4) 
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi8x_xpreheader_bbx_xnphx_xix_xix_xi8_PhiReq/phi_stmt_2847/phi_stmt_2847_sources/type_cast_2850/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi8x_xpreheader_bbx_xnphx_xix_xix_xi8_PhiReq/phi_stmt_2847/phi_stmt_2847_sources/type_cast_2850/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi8x_xpreheader_bbx_xnphx_xix_xix_xi8_PhiReq/phi_stmt_2847/phi_stmt_2847_sources/type_cast_2850/SplitProtocol/Sample/rr
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi8x_xpreheader_bbx_xnphx_xix_xix_xi8_PhiReq/phi_stmt_2847/phi_stmt_2847_sources/type_cast_2850/SplitProtocol/Sample/ra
      -- 
    cp_elements(1728) <= cp_elements(1727);
    -- CP-element group 1729 transition  bypass 
    -- predecessors 1727 
    -- successors 1730 
    -- members (4) 
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi8x_xpreheader_bbx_xnphx_xix_xix_xi8_PhiReq/phi_stmt_2847/phi_stmt_2847_sources/type_cast_2850/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi8x_xpreheader_bbx_xnphx_xix_xix_xi8_PhiReq/phi_stmt_2847/phi_stmt_2847_sources/type_cast_2850/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi8x_xpreheader_bbx_xnphx_xix_xix_xi8_PhiReq/phi_stmt_2847/phi_stmt_2847_sources/type_cast_2850/SplitProtocol/Update/cr
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi8x_xpreheader_bbx_xnphx_xix_xix_xi8_PhiReq/phi_stmt_2847/phi_stmt_2847_sources/type_cast_2850/SplitProtocol/Update/ca
      -- 
    cp_elements(1729) <= cp_elements(1727);
    -- CP-element group 1730 join  transition  bypass 
    -- predecessors 1728 1729 
    -- successors 1737 
    -- members (2) 
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi8x_xpreheader_bbx_xnphx_xix_xix_xi8_PhiReq/phi_stmt_2847/phi_stmt_2847_sources/type_cast_2850/$exit
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi8x_xpreheader_bbx_xnphx_xix_xix_xi8_PhiReq/phi_stmt_2847/phi_stmt_2847_sources/type_cast_2850/SplitProtocol/$exit
      -- 
    cp_element_group_1730: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1730"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1728) & cp_elements(1729);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1730), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1731 fork  transition  bypass 
    -- predecessors 1726 
    -- successors 1732 1734 
    -- members (2) 
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi8x_xpreheader_bbx_xnphx_xix_xix_xi8_PhiReq/phi_stmt_2847/phi_stmt_2847_sources/type_cast_2852/$entry
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi8x_xpreheader_bbx_xnphx_xix_xix_xi8_PhiReq/phi_stmt_2847/phi_stmt_2847_sources/type_cast_2852/SplitProtocol/$entry
      -- 
    cp_elements(1731) <= cp_elements(1726);
    -- CP-element group 1732 transition  output  bypass 
    -- predecessors 1731 
    -- successors 1733 
    -- members (2) 
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi8x_xpreheader_bbx_xnphx_xix_xix_xi8_PhiReq/phi_stmt_2847/phi_stmt_2847_sources/type_cast_2852/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi8x_xpreheader_bbx_xnphx_xix_xix_xi8_PhiReq/phi_stmt_2847/phi_stmt_2847_sources/type_cast_2852/SplitProtocol/Sample/rr
      -- 
    cp_elements(1732) <= cp_elements(1731);
    rr_17403_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1732), ack => type_cast_2852_inst_req_0); -- 
    -- CP-element group 1733 transition  input  bypass 
    -- predecessors 1732 
    -- successors 1736 
    -- members (2) 
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi8x_xpreheader_bbx_xnphx_xix_xix_xi8_PhiReq/phi_stmt_2847/phi_stmt_2847_sources/type_cast_2852/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi8x_xpreheader_bbx_xnphx_xix_xix_xi8_PhiReq/phi_stmt_2847/phi_stmt_2847_sources/type_cast_2852/SplitProtocol/Sample/ra
      -- 
    ra_17404_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2852_inst_ack_0, ack => cp_elements(1733)); -- 
    -- CP-element group 1734 transition  output  bypass 
    -- predecessors 1731 
    -- successors 1735 
    -- members (2) 
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi8x_xpreheader_bbx_xnphx_xix_xix_xi8_PhiReq/phi_stmt_2847/phi_stmt_2847_sources/type_cast_2852/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi8x_xpreheader_bbx_xnphx_xix_xix_xi8_PhiReq/phi_stmt_2847/phi_stmt_2847_sources/type_cast_2852/SplitProtocol/Update/cr
      -- 
    cp_elements(1734) <= cp_elements(1731);
    cr_17408_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1734), ack => type_cast_2852_inst_req_1); -- 
    -- CP-element group 1735 transition  input  bypass 
    -- predecessors 1734 
    -- successors 1736 
    -- members (2) 
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi8x_xpreheader_bbx_xnphx_xix_xix_xi8_PhiReq/phi_stmt_2847/phi_stmt_2847_sources/type_cast_2852/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi8x_xpreheader_bbx_xnphx_xix_xix_xi8_PhiReq/phi_stmt_2847/phi_stmt_2847_sources/type_cast_2852/SplitProtocol/Update/ca
      -- 
    ca_17409_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2852_inst_ack_1, ack => cp_elements(1735)); -- 
    -- CP-element group 1736 join  transition  bypass 
    -- predecessors 1733 1735 
    -- successors 1737 
    -- members (2) 
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi8x_xpreheader_bbx_xnphx_xix_xix_xi8_PhiReq/phi_stmt_2847/phi_stmt_2847_sources/type_cast_2852/$exit
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi8x_xpreheader_bbx_xnphx_xix_xix_xi8_PhiReq/phi_stmt_2847/phi_stmt_2847_sources/type_cast_2852/SplitProtocol/$exit
      -- 
    cp_element_group_1736: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1736"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1733) & cp_elements(1735);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1736), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1737 join  transition  output  bypass 
    -- predecessors 1730 1736 
    -- successors 1742 
    -- members (3) 
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi8x_xpreheader_bbx_xnphx_xix_xix_xi8_PhiReq/phi_stmt_2847/$exit
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi8x_xpreheader_bbx_xnphx_xix_xix_xi8_PhiReq/phi_stmt_2847/phi_stmt_2847_sources/$exit
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi8x_xpreheader_bbx_xnphx_xix_xix_xi8_PhiReq/phi_stmt_2847/phi_stmt_2847_req
      -- 
    cp_element_group_1737: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1737"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1730) & cp_elements(1736);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1737), clk => clk, reset => reset); --
    end block;
    phi_stmt_2847_req_17410_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1737), ack => phi_stmt_2847_req_1); -- 
    -- CP-element group 1738 fork  transition  bypass 
    -- predecessors 1725 
    -- successors 1739 1740 
    -- members (4) 
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi8x_xpreheader_bbx_xnphx_xix_xix_xi8_PhiReq/phi_stmt_2853/$entry
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi8x_xpreheader_bbx_xnphx_xix_xix_xi8_PhiReq/phi_stmt_2853/phi_stmt_2853_sources/$entry
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi8x_xpreheader_bbx_xnphx_xix_xix_xi8_PhiReq/phi_stmt_2853/phi_stmt_2853_sources/type_cast_2856/$entry
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi8x_xpreheader_bbx_xnphx_xix_xix_xi8_PhiReq/phi_stmt_2853/phi_stmt_2853_sources/type_cast_2856/SplitProtocol/$entry
      -- 
    cp_elements(1738) <= cp_elements(1725);
    -- CP-element group 1739 transition  bypass 
    -- predecessors 1738 
    -- successors 1741 
    -- members (4) 
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi8x_xpreheader_bbx_xnphx_xix_xix_xi8_PhiReq/phi_stmt_2853/phi_stmt_2853_sources/type_cast_2856/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi8x_xpreheader_bbx_xnphx_xix_xix_xi8_PhiReq/phi_stmt_2853/phi_stmt_2853_sources/type_cast_2856/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi8x_xpreheader_bbx_xnphx_xix_xix_xi8_PhiReq/phi_stmt_2853/phi_stmt_2853_sources/type_cast_2856/SplitProtocol/Sample/rr
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi8x_xpreheader_bbx_xnphx_xix_xix_xi8_PhiReq/phi_stmt_2853/phi_stmt_2853_sources/type_cast_2856/SplitProtocol/Sample/ra
      -- 
    cp_elements(1739) <= cp_elements(1738);
    -- CP-element group 1740 transition  bypass 
    -- predecessors 1738 
    -- successors 1741 
    -- members (4) 
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi8x_xpreheader_bbx_xnphx_xix_xix_xi8_PhiReq/phi_stmt_2853/phi_stmt_2853_sources/type_cast_2856/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi8x_xpreheader_bbx_xnphx_xix_xix_xi8_PhiReq/phi_stmt_2853/phi_stmt_2853_sources/type_cast_2856/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi8x_xpreheader_bbx_xnphx_xix_xix_xi8_PhiReq/phi_stmt_2853/phi_stmt_2853_sources/type_cast_2856/SplitProtocol/Update/cr
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi8x_xpreheader_bbx_xnphx_xix_xix_xi8_PhiReq/phi_stmt_2853/phi_stmt_2853_sources/type_cast_2856/SplitProtocol/Update/ca
      -- 
    cp_elements(1740) <= cp_elements(1738);
    -- CP-element group 1741 join  transition  output  bypass 
    -- predecessors 1739 1740 
    -- successors 1742 
    -- members (5) 
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi8x_xpreheader_bbx_xnphx_xix_xix_xi8_PhiReq/phi_stmt_2853/$exit
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi8x_xpreheader_bbx_xnphx_xix_xix_xi8_PhiReq/phi_stmt_2853/phi_stmt_2853_sources/$exit
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi8x_xpreheader_bbx_xnphx_xix_xix_xi8_PhiReq/phi_stmt_2853/phi_stmt_2853_sources/type_cast_2856/$exit
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi8x_xpreheader_bbx_xnphx_xix_xix_xi8_PhiReq/phi_stmt_2853/phi_stmt_2853_sources/type_cast_2856/SplitProtocol/$exit
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi8x_xpreheader_bbx_xnphx_xix_xix_xi8_PhiReq/phi_stmt_2853/phi_stmt_2853_req
      -- 
    cp_element_group_1741: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1741"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1739) & cp_elements(1740);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1741), clk => clk, reset => reset); --
    end block;
    phi_stmt_2853_req_17433_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1741), ack => phi_stmt_2853_req_1); -- 
    -- CP-element group 1742 join  transition  bypass 
    -- predecessors 1737 1741 
    -- successors 1743 
    -- members (1) 
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi8x_xpreheader_bbx_xnphx_xix_xix_xi8_PhiReq/$exit
      -- 
    cp_element_group_1742: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1742"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1737) & cp_elements(1741);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1742), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1743 merge  place  bypass 
    -- predecessors 1724 1742 
    -- successors 1744 
    -- members (1) 
      -- 	branch_block_stmt_2042/merge_stmt_2846_PhiReqMerge
      -- 
    cp_elements(1743) <= OrReduce(cp_elements(1724) & cp_elements(1742));
    -- CP-element group 1744 fork  transition  bypass 
    -- predecessors 1743 
    -- successors 1745 1746 
    -- members (1) 
      -- 	branch_block_stmt_2042/merge_stmt_2846_PhiAck/$entry
      -- 
    cp_elements(1744) <= cp_elements(1743);
    -- CP-element group 1745 transition  input  bypass 
    -- predecessors 1744 
    -- successors 1747 
    -- members (1) 
      -- 	branch_block_stmt_2042/merge_stmt_2846_PhiAck/phi_stmt_2847_ack
      -- 
    phi_stmt_2847_ack_17438_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2847_ack_0, ack => cp_elements(1745)); -- 
    -- CP-element group 1746 transition  input  bypass 
    -- predecessors 1744 
    -- successors 1747 
    -- members (1) 
      -- 	branch_block_stmt_2042/merge_stmt_2846_PhiAck/phi_stmt_2853_ack
      -- 
    phi_stmt_2853_ack_17439_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2853_ack_0, ack => cp_elements(1746)); -- 
    -- CP-element group 1747 join  transition  bypass 
    -- predecessors 1745 1746 
    -- successors 32 
    -- members (1) 
      -- 	branch_block_stmt_2042/merge_stmt_2846_PhiAck/$exit
      -- 
    cp_element_group_1747: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1747"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1745) & cp_elements(1746);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1747), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1748 fork  transition  bypass 
    -- predecessors 598 
    -- successors 1749 1755 
    -- members (1) 
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi8_xx_x_crit_edgex_xix_xix_xi11x_xloopexit_PhiReq/$entry
      -- 
    cp_elements(1748) <= cp_elements(598);
    -- CP-element group 1749 fork  transition  bypass 
    -- predecessors 1748 
    -- successors 1750 1752 
    -- members (4) 
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi8_xx_x_crit_edgex_xix_xix_xi11x_xloopexit_PhiReq/phi_stmt_2885/$entry
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi8_xx_x_crit_edgex_xix_xix_xi11x_xloopexit_PhiReq/phi_stmt_2885/phi_stmt_2885_sources/$entry
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi8_xx_x_crit_edgex_xix_xix_xi11x_xloopexit_PhiReq/phi_stmt_2885/phi_stmt_2885_sources/type_cast_2888/$entry
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi8_xx_x_crit_edgex_xix_xix_xi11x_xloopexit_PhiReq/phi_stmt_2885/phi_stmt_2885_sources/type_cast_2888/SplitProtocol/$entry
      -- 
    cp_elements(1749) <= cp_elements(1748);
    -- CP-element group 1750 transition  output  bypass 
    -- predecessors 1749 
    -- successors 1751 
    -- members (2) 
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi8_xx_x_crit_edgex_xix_xix_xi11x_xloopexit_PhiReq/phi_stmt_2885/phi_stmt_2885_sources/type_cast_2888/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi8_xx_x_crit_edgex_xix_xix_xi11x_xloopexit_PhiReq/phi_stmt_2885/phi_stmt_2885_sources/type_cast_2888/SplitProtocol/Sample/rr
      -- 
    cp_elements(1750) <= cp_elements(1749);
    rr_17462_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1750), ack => type_cast_2888_inst_req_0); -- 
    -- CP-element group 1751 transition  input  bypass 
    -- predecessors 1750 
    -- successors 1754 
    -- members (2) 
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi8_xx_x_crit_edgex_xix_xix_xi11x_xloopexit_PhiReq/phi_stmt_2885/phi_stmt_2885_sources/type_cast_2888/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi8_xx_x_crit_edgex_xix_xix_xi11x_xloopexit_PhiReq/phi_stmt_2885/phi_stmt_2885_sources/type_cast_2888/SplitProtocol/Sample/ra
      -- 
    ra_17463_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2888_inst_ack_0, ack => cp_elements(1751)); -- 
    -- CP-element group 1752 transition  output  bypass 
    -- predecessors 1749 
    -- successors 1753 
    -- members (2) 
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi8_xx_x_crit_edgex_xix_xix_xi11x_xloopexit_PhiReq/phi_stmt_2885/phi_stmt_2885_sources/type_cast_2888/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi8_xx_x_crit_edgex_xix_xix_xi11x_xloopexit_PhiReq/phi_stmt_2885/phi_stmt_2885_sources/type_cast_2888/SplitProtocol/Update/cr
      -- 
    cp_elements(1752) <= cp_elements(1749);
    cr_17467_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1752), ack => type_cast_2888_inst_req_1); -- 
    -- CP-element group 1753 transition  input  bypass 
    -- predecessors 1752 
    -- successors 1754 
    -- members (2) 
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi8_xx_x_crit_edgex_xix_xix_xi11x_xloopexit_PhiReq/phi_stmt_2885/phi_stmt_2885_sources/type_cast_2888/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi8_xx_x_crit_edgex_xix_xix_xi11x_xloopexit_PhiReq/phi_stmt_2885/phi_stmt_2885_sources/type_cast_2888/SplitProtocol/Update/ca
      -- 
    ca_17468_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2888_inst_ack_1, ack => cp_elements(1753)); -- 
    -- CP-element group 1754 join  transition  output  bypass 
    -- predecessors 1751 1753 
    -- successors 1761 
    -- members (5) 
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi8_xx_x_crit_edgex_xix_xix_xi11x_xloopexit_PhiReq/phi_stmt_2885/$exit
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi8_xx_x_crit_edgex_xix_xix_xi11x_xloopexit_PhiReq/phi_stmt_2885/phi_stmt_2885_sources/$exit
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi8_xx_x_crit_edgex_xix_xix_xi11x_xloopexit_PhiReq/phi_stmt_2885/phi_stmt_2885_sources/type_cast_2888/$exit
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi8_xx_x_crit_edgex_xix_xix_xi11x_xloopexit_PhiReq/phi_stmt_2885/phi_stmt_2885_sources/type_cast_2888/SplitProtocol/$exit
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi8_xx_x_crit_edgex_xix_xix_xi11x_xloopexit_PhiReq/phi_stmt_2885/phi_stmt_2885_req
      -- 
    cp_element_group_1754: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1754"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1751) & cp_elements(1753);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1754), clk => clk, reset => reset); --
    end block;
    phi_stmt_2885_req_17469_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1754), ack => phi_stmt_2885_req_0); -- 
    -- CP-element group 1755 fork  transition  bypass 
    -- predecessors 1748 
    -- successors 1756 1758 
    -- members (4) 
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi8_xx_x_crit_edgex_xix_xix_xi11x_xloopexit_PhiReq/phi_stmt_2889/$entry
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi8_xx_x_crit_edgex_xix_xix_xi11x_xloopexit_PhiReq/phi_stmt_2889/phi_stmt_2889_sources/$entry
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi8_xx_x_crit_edgex_xix_xix_xi11x_xloopexit_PhiReq/phi_stmt_2889/phi_stmt_2889_sources/type_cast_2892/$entry
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi8_xx_x_crit_edgex_xix_xix_xi11x_xloopexit_PhiReq/phi_stmt_2889/phi_stmt_2889_sources/type_cast_2892/SplitProtocol/$entry
      -- 
    cp_elements(1755) <= cp_elements(1748);
    -- CP-element group 1756 transition  output  bypass 
    -- predecessors 1755 
    -- successors 1757 
    -- members (2) 
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi8_xx_x_crit_edgex_xix_xix_xi11x_xloopexit_PhiReq/phi_stmt_2889/phi_stmt_2889_sources/type_cast_2892/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi8_xx_x_crit_edgex_xix_xix_xi11x_xloopexit_PhiReq/phi_stmt_2889/phi_stmt_2889_sources/type_cast_2892/SplitProtocol/Sample/rr
      -- 
    cp_elements(1756) <= cp_elements(1755);
    rr_17485_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1756), ack => type_cast_2892_inst_req_0); -- 
    -- CP-element group 1757 transition  input  bypass 
    -- predecessors 1756 
    -- successors 1760 
    -- members (2) 
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi8_xx_x_crit_edgex_xix_xix_xi11x_xloopexit_PhiReq/phi_stmt_2889/phi_stmt_2889_sources/type_cast_2892/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi8_xx_x_crit_edgex_xix_xix_xi11x_xloopexit_PhiReq/phi_stmt_2889/phi_stmt_2889_sources/type_cast_2892/SplitProtocol/Sample/ra
      -- 
    ra_17486_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2892_inst_ack_0, ack => cp_elements(1757)); -- 
    -- CP-element group 1758 transition  output  bypass 
    -- predecessors 1755 
    -- successors 1759 
    -- members (2) 
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi8_xx_x_crit_edgex_xix_xix_xi11x_xloopexit_PhiReq/phi_stmt_2889/phi_stmt_2889_sources/type_cast_2892/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi8_xx_x_crit_edgex_xix_xix_xi11x_xloopexit_PhiReq/phi_stmt_2889/phi_stmt_2889_sources/type_cast_2892/SplitProtocol/Update/cr
      -- 
    cp_elements(1758) <= cp_elements(1755);
    cr_17490_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1758), ack => type_cast_2892_inst_req_1); -- 
    -- CP-element group 1759 transition  input  bypass 
    -- predecessors 1758 
    -- successors 1760 
    -- members (2) 
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi8_xx_x_crit_edgex_xix_xix_xi11x_xloopexit_PhiReq/phi_stmt_2889/phi_stmt_2889_sources/type_cast_2892/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi8_xx_x_crit_edgex_xix_xix_xi11x_xloopexit_PhiReq/phi_stmt_2889/phi_stmt_2889_sources/type_cast_2892/SplitProtocol/Update/ca
      -- 
    ca_17491_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2892_inst_ack_1, ack => cp_elements(1759)); -- 
    -- CP-element group 1760 join  transition  output  bypass 
    -- predecessors 1757 1759 
    -- successors 1761 
    -- members (5) 
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi8_xx_x_crit_edgex_xix_xix_xi11x_xloopexit_PhiReq/phi_stmt_2889/$exit
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi8_xx_x_crit_edgex_xix_xix_xi11x_xloopexit_PhiReq/phi_stmt_2889/phi_stmt_2889_sources/$exit
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi8_xx_x_crit_edgex_xix_xix_xi11x_xloopexit_PhiReq/phi_stmt_2889/phi_stmt_2889_sources/type_cast_2892/$exit
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi8_xx_x_crit_edgex_xix_xix_xi11x_xloopexit_PhiReq/phi_stmt_2889/phi_stmt_2889_sources/type_cast_2892/SplitProtocol/$exit
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi8_xx_x_crit_edgex_xix_xix_xi11x_xloopexit_PhiReq/phi_stmt_2889/phi_stmt_2889_req
      -- 
    cp_element_group_1760: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1760"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1757) & cp_elements(1759);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1760), clk => clk, reset => reset); --
    end block;
    phi_stmt_2889_req_17492_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1760), ack => phi_stmt_2889_req_0); -- 
    -- CP-element group 1761 join  transition  bypass 
    -- predecessors 1754 1760 
    -- successors 1762 
    -- members (1) 
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi8_xx_x_crit_edgex_xix_xix_xi11x_xloopexit_PhiReq/$exit
      -- 
    cp_element_group_1761: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1761"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1754) & cp_elements(1760);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1761), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1762 place  bypass 
    -- predecessors 1761 
    -- successors 1763 
    -- members (1) 
      -- 	branch_block_stmt_2042/merge_stmt_2884_PhiReqMerge
      -- 
    cp_elements(1762) <= cp_elements(1761);
    -- CP-element group 1763 fork  transition  bypass 
    -- predecessors 1762 
    -- successors 1764 1765 
    -- members (1) 
      -- 	branch_block_stmt_2042/merge_stmt_2884_PhiAck/$entry
      -- 
    cp_elements(1763) <= cp_elements(1762);
    -- CP-element group 1764 transition  input  bypass 
    -- predecessors 1763 
    -- successors 1766 
    -- members (1) 
      -- 	branch_block_stmt_2042/merge_stmt_2884_PhiAck/phi_stmt_2885_ack
      -- 
    phi_stmt_2885_ack_17497_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2885_ack_0, ack => cp_elements(1764)); -- 
    -- CP-element group 1765 transition  input  bypass 
    -- predecessors 1763 
    -- successors 1766 
    -- members (1) 
      -- 	branch_block_stmt_2042/merge_stmt_2884_PhiAck/phi_stmt_2889_ack
      -- 
    phi_stmt_2889_ack_17498_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2889_ack_0, ack => cp_elements(1765)); -- 
    -- CP-element group 1766 join  transition  bypass 
    -- predecessors 1764 1765 
    -- successors 34 
    -- members (1) 
      -- 	branch_block_stmt_2042/merge_stmt_2884_PhiAck/$exit
      -- 
    cp_element_group_1766: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1766"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1764) & cp_elements(1765);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1766), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1767 fork  transition  bypass 
    -- predecessors 576 
    -- successors 1768 1780 
    -- members (1) 
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xix_xi5_xx_x_crit_edgex_xix_xix_xi11_PhiReq/$entry
      -- 
    cp_elements(1767) <= cp_elements(576);
    -- CP-element group 1768 fork  transition  bypass 
    -- predecessors 1767 
    -- successors 1769 1775 
    -- members (2) 
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xix_xi5_xx_x_crit_edgex_xix_xix_xi11_PhiReq/phi_stmt_2896/$entry
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xix_xi5_xx_x_crit_edgex_xix_xix_xi11_PhiReq/phi_stmt_2896/phi_stmt_2896_sources/$entry
      -- 
    cp_elements(1768) <= cp_elements(1767);
    -- CP-element group 1769 fork  transition  bypass 
    -- predecessors 1768 
    -- successors 1770 1772 
    -- members (2) 
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xix_xi5_xx_x_crit_edgex_xix_xix_xi11_PhiReq/phi_stmt_2896/phi_stmt_2896_sources/type_cast_2899/$entry
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xix_xi5_xx_x_crit_edgex_xix_xix_xi11_PhiReq/phi_stmt_2896/phi_stmt_2896_sources/type_cast_2899/SplitProtocol/$entry
      -- 
    cp_elements(1769) <= cp_elements(1768);
    -- CP-element group 1770 transition  output  bypass 
    -- predecessors 1769 
    -- successors 1771 
    -- members (2) 
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xix_xi5_xx_x_crit_edgex_xix_xix_xi11_PhiReq/phi_stmt_2896/phi_stmt_2896_sources/type_cast_2899/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xix_xi5_xx_x_crit_edgex_xix_xix_xi11_PhiReq/phi_stmt_2896/phi_stmt_2896_sources/type_cast_2899/SplitProtocol/Sample/rr
      -- 
    cp_elements(1770) <= cp_elements(1769);
    rr_17517_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1770), ack => type_cast_2899_inst_req_0); -- 
    -- CP-element group 1771 transition  input  bypass 
    -- predecessors 1770 
    -- successors 1774 
    -- members (2) 
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xix_xi5_xx_x_crit_edgex_xix_xix_xi11_PhiReq/phi_stmt_2896/phi_stmt_2896_sources/type_cast_2899/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xix_xi5_xx_x_crit_edgex_xix_xix_xi11_PhiReq/phi_stmt_2896/phi_stmt_2896_sources/type_cast_2899/SplitProtocol/Sample/ra
      -- 
    ra_17518_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2899_inst_ack_0, ack => cp_elements(1771)); -- 
    -- CP-element group 1772 transition  output  bypass 
    -- predecessors 1769 
    -- successors 1773 
    -- members (2) 
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xix_xi5_xx_x_crit_edgex_xix_xix_xi11_PhiReq/phi_stmt_2896/phi_stmt_2896_sources/type_cast_2899/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xix_xi5_xx_x_crit_edgex_xix_xix_xi11_PhiReq/phi_stmt_2896/phi_stmt_2896_sources/type_cast_2899/SplitProtocol/Update/cr
      -- 
    cp_elements(1772) <= cp_elements(1769);
    cr_17522_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1772), ack => type_cast_2899_inst_req_1); -- 
    -- CP-element group 1773 transition  input  bypass 
    -- predecessors 1772 
    -- successors 1774 
    -- members (2) 
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xix_xi5_xx_x_crit_edgex_xix_xix_xi11_PhiReq/phi_stmt_2896/phi_stmt_2896_sources/type_cast_2899/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xix_xi5_xx_x_crit_edgex_xix_xix_xi11_PhiReq/phi_stmt_2896/phi_stmt_2896_sources/type_cast_2899/SplitProtocol/Update/ca
      -- 
    ca_17523_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2899_inst_ack_1, ack => cp_elements(1773)); -- 
    -- CP-element group 1774 join  transition  bypass 
    -- predecessors 1771 1773 
    -- successors 1779 
    -- members (2) 
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xix_xi5_xx_x_crit_edgex_xix_xix_xi11_PhiReq/phi_stmt_2896/phi_stmt_2896_sources/type_cast_2899/$exit
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xix_xi5_xx_x_crit_edgex_xix_xix_xi11_PhiReq/phi_stmt_2896/phi_stmt_2896_sources/type_cast_2899/SplitProtocol/$exit
      -- 
    cp_element_group_1774: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1774"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1771) & cp_elements(1773);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1774), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1775 fork  transition  bypass 
    -- predecessors 1768 
    -- successors 1776 1777 
    -- members (2) 
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xix_xi5_xx_x_crit_edgex_xix_xix_xi11_PhiReq/phi_stmt_2896/phi_stmt_2896_sources/type_cast_2901/$entry
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xix_xi5_xx_x_crit_edgex_xix_xix_xi11_PhiReq/phi_stmt_2896/phi_stmt_2896_sources/type_cast_2901/SplitProtocol/$entry
      -- 
    cp_elements(1775) <= cp_elements(1768);
    -- CP-element group 1776 transition  bypass 
    -- predecessors 1775 
    -- successors 1778 
    -- members (4) 
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xix_xi5_xx_x_crit_edgex_xix_xix_xi11_PhiReq/phi_stmt_2896/phi_stmt_2896_sources/type_cast_2901/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xix_xi5_xx_x_crit_edgex_xix_xix_xi11_PhiReq/phi_stmt_2896/phi_stmt_2896_sources/type_cast_2901/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xix_xi5_xx_x_crit_edgex_xix_xix_xi11_PhiReq/phi_stmt_2896/phi_stmt_2896_sources/type_cast_2901/SplitProtocol/Sample/rr
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xix_xi5_xx_x_crit_edgex_xix_xix_xi11_PhiReq/phi_stmt_2896/phi_stmt_2896_sources/type_cast_2901/SplitProtocol/Sample/ra
      -- 
    cp_elements(1776) <= cp_elements(1775);
    -- CP-element group 1777 transition  bypass 
    -- predecessors 1775 
    -- successors 1778 
    -- members (4) 
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xix_xi5_xx_x_crit_edgex_xix_xix_xi11_PhiReq/phi_stmt_2896/phi_stmt_2896_sources/type_cast_2901/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xix_xi5_xx_x_crit_edgex_xix_xix_xi11_PhiReq/phi_stmt_2896/phi_stmt_2896_sources/type_cast_2901/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xix_xi5_xx_x_crit_edgex_xix_xix_xi11_PhiReq/phi_stmt_2896/phi_stmt_2896_sources/type_cast_2901/SplitProtocol/Update/cr
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xix_xi5_xx_x_crit_edgex_xix_xix_xi11_PhiReq/phi_stmt_2896/phi_stmt_2896_sources/type_cast_2901/SplitProtocol/Update/ca
      -- 
    cp_elements(1777) <= cp_elements(1775);
    -- CP-element group 1778 join  transition  bypass 
    -- predecessors 1776 1777 
    -- successors 1779 
    -- members (2) 
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xix_xi5_xx_x_crit_edgex_xix_xix_xi11_PhiReq/phi_stmt_2896/phi_stmt_2896_sources/type_cast_2901/$exit
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xix_xi5_xx_x_crit_edgex_xix_xix_xi11_PhiReq/phi_stmt_2896/phi_stmt_2896_sources/type_cast_2901/SplitProtocol/$exit
      -- 
    cp_element_group_1778: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1778"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1776) & cp_elements(1777);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1778), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1779 join  transition  output  bypass 
    -- predecessors 1774 1778 
    -- successors 1784 
    -- members (3) 
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xix_xi5_xx_x_crit_edgex_xix_xix_xi11_PhiReq/phi_stmt_2896/$exit
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xix_xi5_xx_x_crit_edgex_xix_xix_xi11_PhiReq/phi_stmt_2896/phi_stmt_2896_sources/$exit
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xix_xi5_xx_x_crit_edgex_xix_xix_xi11_PhiReq/phi_stmt_2896/phi_stmt_2896_req
      -- 
    cp_element_group_1779: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1779"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1774) & cp_elements(1778);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1779), clk => clk, reset => reset); --
    end block;
    phi_stmt_2896_req_17540_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1779), ack => phi_stmt_2896_req_0); -- 
    -- CP-element group 1780 fork  transition  bypass 
    -- predecessors 1767 
    -- successors 1781 1782 
    -- members (4) 
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xix_xi5_xx_x_crit_edgex_xix_xix_xi11_PhiReq/phi_stmt_2902/$entry
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xix_xi5_xx_x_crit_edgex_xix_xix_xi11_PhiReq/phi_stmt_2902/phi_stmt_2902_sources/$entry
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xix_xi5_xx_x_crit_edgex_xix_xix_xi11_PhiReq/phi_stmt_2902/phi_stmt_2902_sources/type_cast_2908/$entry
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xix_xi5_xx_x_crit_edgex_xix_xix_xi11_PhiReq/phi_stmt_2902/phi_stmt_2902_sources/type_cast_2908/SplitProtocol/$entry
      -- 
    cp_elements(1780) <= cp_elements(1767);
    -- CP-element group 1781 transition  bypass 
    -- predecessors 1780 
    -- successors 1783 
    -- members (4) 
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xix_xi5_xx_x_crit_edgex_xix_xix_xi11_PhiReq/phi_stmt_2902/phi_stmt_2902_sources/type_cast_2908/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xix_xi5_xx_x_crit_edgex_xix_xix_xi11_PhiReq/phi_stmt_2902/phi_stmt_2902_sources/type_cast_2908/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xix_xi5_xx_x_crit_edgex_xix_xix_xi11_PhiReq/phi_stmt_2902/phi_stmt_2902_sources/type_cast_2908/SplitProtocol/Sample/rr
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xix_xi5_xx_x_crit_edgex_xix_xix_xi11_PhiReq/phi_stmt_2902/phi_stmt_2902_sources/type_cast_2908/SplitProtocol/Sample/ra
      -- 
    cp_elements(1781) <= cp_elements(1780);
    -- CP-element group 1782 transition  bypass 
    -- predecessors 1780 
    -- successors 1783 
    -- members (4) 
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xix_xi5_xx_x_crit_edgex_xix_xix_xi11_PhiReq/phi_stmt_2902/phi_stmt_2902_sources/type_cast_2908/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xix_xi5_xx_x_crit_edgex_xix_xix_xi11_PhiReq/phi_stmt_2902/phi_stmt_2902_sources/type_cast_2908/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xix_xi5_xx_x_crit_edgex_xix_xix_xi11_PhiReq/phi_stmt_2902/phi_stmt_2902_sources/type_cast_2908/SplitProtocol/Update/cr
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xix_xi5_xx_x_crit_edgex_xix_xix_xi11_PhiReq/phi_stmt_2902/phi_stmt_2902_sources/type_cast_2908/SplitProtocol/Update/ca
      -- 
    cp_elements(1782) <= cp_elements(1780);
    -- CP-element group 1783 join  transition  output  bypass 
    -- predecessors 1781 1782 
    -- successors 1784 
    -- members (5) 
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xix_xi5_xx_x_crit_edgex_xix_xix_xi11_PhiReq/phi_stmt_2902/$exit
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xix_xi5_xx_x_crit_edgex_xix_xix_xi11_PhiReq/phi_stmt_2902/phi_stmt_2902_sources/$exit
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xix_xi5_xx_x_crit_edgex_xix_xix_xi11_PhiReq/phi_stmt_2902/phi_stmt_2902_sources/type_cast_2908/$exit
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xix_xi5_xx_x_crit_edgex_xix_xix_xi11_PhiReq/phi_stmt_2902/phi_stmt_2902_sources/type_cast_2908/SplitProtocol/$exit
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xix_xi5_xx_x_crit_edgex_xix_xix_xi11_PhiReq/phi_stmt_2902/phi_stmt_2902_req
      -- 
    cp_element_group_1783: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1783"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1781) & cp_elements(1782);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1783), clk => clk, reset => reset); --
    end block;
    phi_stmt_2902_req_17563_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1783), ack => phi_stmt_2902_req_0); -- 
    -- CP-element group 1784 join  transition  bypass 
    -- predecessors 1779 1783 
    -- successors 1805 
    -- members (1) 
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xix_xi5_xx_x_crit_edgex_xix_xix_xi11_PhiReq/$exit
      -- 
    cp_element_group_1784: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1784"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1779) & cp_elements(1783);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1784), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1785 fork  transition  bypass 
    -- predecessors 34 
    -- successors 1786 1798 
    -- members (1) 
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi11x_xloopexit_xx_x_crit_edgex_xix_xix_xi11_PhiReq/$entry
      -- 
    cp_elements(1785) <= cp_elements(34);
    -- CP-element group 1786 fork  transition  bypass 
    -- predecessors 1785 
    -- successors 1787 1791 
    -- members (2) 
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi11x_xloopexit_xx_x_crit_edgex_xix_xix_xi11_PhiReq/phi_stmt_2896/$entry
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi11x_xloopexit_xx_x_crit_edgex_xix_xix_xi11_PhiReq/phi_stmt_2896/phi_stmt_2896_sources/$entry
      -- 
    cp_elements(1786) <= cp_elements(1785);
    -- CP-element group 1787 fork  transition  bypass 
    -- predecessors 1786 
    -- successors 1788 1789 
    -- members (2) 
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi11x_xloopexit_xx_x_crit_edgex_xix_xix_xi11_PhiReq/phi_stmt_2896/phi_stmt_2896_sources/type_cast_2899/$entry
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi11x_xloopexit_xx_x_crit_edgex_xix_xix_xi11_PhiReq/phi_stmt_2896/phi_stmt_2896_sources/type_cast_2899/SplitProtocol/$entry
      -- 
    cp_elements(1787) <= cp_elements(1786);
    -- CP-element group 1788 transition  bypass 
    -- predecessors 1787 
    -- successors 1790 
    -- members (4) 
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi11x_xloopexit_xx_x_crit_edgex_xix_xix_xi11_PhiReq/phi_stmt_2896/phi_stmt_2896_sources/type_cast_2899/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi11x_xloopexit_xx_x_crit_edgex_xix_xix_xi11_PhiReq/phi_stmt_2896/phi_stmt_2896_sources/type_cast_2899/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi11x_xloopexit_xx_x_crit_edgex_xix_xix_xi11_PhiReq/phi_stmt_2896/phi_stmt_2896_sources/type_cast_2899/SplitProtocol/Sample/rr
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi11x_xloopexit_xx_x_crit_edgex_xix_xix_xi11_PhiReq/phi_stmt_2896/phi_stmt_2896_sources/type_cast_2899/SplitProtocol/Sample/ra
      -- 
    cp_elements(1788) <= cp_elements(1787);
    -- CP-element group 1789 transition  bypass 
    -- predecessors 1787 
    -- successors 1790 
    -- members (4) 
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi11x_xloopexit_xx_x_crit_edgex_xix_xix_xi11_PhiReq/phi_stmt_2896/phi_stmt_2896_sources/type_cast_2899/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi11x_xloopexit_xx_x_crit_edgex_xix_xix_xi11_PhiReq/phi_stmt_2896/phi_stmt_2896_sources/type_cast_2899/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi11x_xloopexit_xx_x_crit_edgex_xix_xix_xi11_PhiReq/phi_stmt_2896/phi_stmt_2896_sources/type_cast_2899/SplitProtocol/Update/cr
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi11x_xloopexit_xx_x_crit_edgex_xix_xix_xi11_PhiReq/phi_stmt_2896/phi_stmt_2896_sources/type_cast_2899/SplitProtocol/Update/ca
      -- 
    cp_elements(1789) <= cp_elements(1787);
    -- CP-element group 1790 join  transition  bypass 
    -- predecessors 1788 1789 
    -- successors 1797 
    -- members (2) 
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi11x_xloopexit_xx_x_crit_edgex_xix_xix_xi11_PhiReq/phi_stmt_2896/phi_stmt_2896_sources/type_cast_2899/$exit
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi11x_xloopexit_xx_x_crit_edgex_xix_xix_xi11_PhiReq/phi_stmt_2896/phi_stmt_2896_sources/type_cast_2899/SplitProtocol/$exit
      -- 
    cp_element_group_1790: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1790"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1788) & cp_elements(1789);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1790), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1791 fork  transition  bypass 
    -- predecessors 1786 
    -- successors 1792 1794 
    -- members (2) 
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi11x_xloopexit_xx_x_crit_edgex_xix_xix_xi11_PhiReq/phi_stmt_2896/phi_stmt_2896_sources/type_cast_2901/$entry
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi11x_xloopexit_xx_x_crit_edgex_xix_xix_xi11_PhiReq/phi_stmt_2896/phi_stmt_2896_sources/type_cast_2901/SplitProtocol/$entry
      -- 
    cp_elements(1791) <= cp_elements(1786);
    -- CP-element group 1792 transition  output  bypass 
    -- predecessors 1791 
    -- successors 1793 
    -- members (2) 
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi11x_xloopexit_xx_x_crit_edgex_xix_xix_xi11_PhiReq/phi_stmt_2896/phi_stmt_2896_sources/type_cast_2901/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi11x_xloopexit_xx_x_crit_edgex_xix_xix_xi11_PhiReq/phi_stmt_2896/phi_stmt_2896_sources/type_cast_2901/SplitProtocol/Sample/rr
      -- 
    cp_elements(1792) <= cp_elements(1791);
    rr_17598_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1792), ack => type_cast_2901_inst_req_0); -- 
    -- CP-element group 1793 transition  input  bypass 
    -- predecessors 1792 
    -- successors 1796 
    -- members (2) 
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi11x_xloopexit_xx_x_crit_edgex_xix_xix_xi11_PhiReq/phi_stmt_2896/phi_stmt_2896_sources/type_cast_2901/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi11x_xloopexit_xx_x_crit_edgex_xix_xix_xi11_PhiReq/phi_stmt_2896/phi_stmt_2896_sources/type_cast_2901/SplitProtocol/Sample/ra
      -- 
    ra_17599_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2901_inst_ack_0, ack => cp_elements(1793)); -- 
    -- CP-element group 1794 transition  output  bypass 
    -- predecessors 1791 
    -- successors 1795 
    -- members (2) 
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi11x_xloopexit_xx_x_crit_edgex_xix_xix_xi11_PhiReq/phi_stmt_2896/phi_stmt_2896_sources/type_cast_2901/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi11x_xloopexit_xx_x_crit_edgex_xix_xix_xi11_PhiReq/phi_stmt_2896/phi_stmt_2896_sources/type_cast_2901/SplitProtocol/Update/cr
      -- 
    cp_elements(1794) <= cp_elements(1791);
    cr_17603_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1794), ack => type_cast_2901_inst_req_1); -- 
    -- CP-element group 1795 transition  input  bypass 
    -- predecessors 1794 
    -- successors 1796 
    -- members (2) 
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi11x_xloopexit_xx_x_crit_edgex_xix_xix_xi11_PhiReq/phi_stmt_2896/phi_stmt_2896_sources/type_cast_2901/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi11x_xloopexit_xx_x_crit_edgex_xix_xix_xi11_PhiReq/phi_stmt_2896/phi_stmt_2896_sources/type_cast_2901/SplitProtocol/Update/ca
      -- 
    ca_17604_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2901_inst_ack_1, ack => cp_elements(1795)); -- 
    -- CP-element group 1796 join  transition  bypass 
    -- predecessors 1793 1795 
    -- successors 1797 
    -- members (2) 
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi11x_xloopexit_xx_x_crit_edgex_xix_xix_xi11_PhiReq/phi_stmt_2896/phi_stmt_2896_sources/type_cast_2901/$exit
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi11x_xloopexit_xx_x_crit_edgex_xix_xix_xi11_PhiReq/phi_stmt_2896/phi_stmt_2896_sources/type_cast_2901/SplitProtocol/$exit
      -- 
    cp_element_group_1796: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1796"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1793) & cp_elements(1795);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1796), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1797 join  transition  output  bypass 
    -- predecessors 1790 1796 
    -- successors 1804 
    -- members (3) 
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi11x_xloopexit_xx_x_crit_edgex_xix_xix_xi11_PhiReq/phi_stmt_2896/$exit
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi11x_xloopexit_xx_x_crit_edgex_xix_xix_xi11_PhiReq/phi_stmt_2896/phi_stmt_2896_sources/$exit
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi11x_xloopexit_xx_x_crit_edgex_xix_xix_xi11_PhiReq/phi_stmt_2896/phi_stmt_2896_req
      -- 
    cp_element_group_1797: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1797"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1790) & cp_elements(1796);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1797), clk => clk, reset => reset); --
    end block;
    phi_stmt_2896_req_17605_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1797), ack => phi_stmt_2896_req_1); -- 
    -- CP-element group 1798 fork  transition  bypass 
    -- predecessors 1785 
    -- successors 1799 1801 
    -- members (4) 
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi11x_xloopexit_xx_x_crit_edgex_xix_xix_xi11_PhiReq/phi_stmt_2902/$entry
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi11x_xloopexit_xx_x_crit_edgex_xix_xix_xi11_PhiReq/phi_stmt_2902/phi_stmt_2902_sources/$entry
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi11x_xloopexit_xx_x_crit_edgex_xix_xix_xi11_PhiReq/phi_stmt_2902/phi_stmt_2902_sources/type_cast_2908/$entry
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi11x_xloopexit_xx_x_crit_edgex_xix_xix_xi11_PhiReq/phi_stmt_2902/phi_stmt_2902_sources/type_cast_2908/SplitProtocol/$entry
      -- 
    cp_elements(1798) <= cp_elements(1785);
    -- CP-element group 1799 transition  output  bypass 
    -- predecessors 1798 
    -- successors 1800 
    -- members (2) 
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi11x_xloopexit_xx_x_crit_edgex_xix_xix_xi11_PhiReq/phi_stmt_2902/phi_stmt_2902_sources/type_cast_2908/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi11x_xloopexit_xx_x_crit_edgex_xix_xix_xi11_PhiReq/phi_stmt_2902/phi_stmt_2902_sources/type_cast_2908/SplitProtocol/Sample/rr
      -- 
    cp_elements(1799) <= cp_elements(1798);
    rr_17621_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1799), ack => type_cast_2908_inst_req_0); -- 
    -- CP-element group 1800 transition  input  bypass 
    -- predecessors 1799 
    -- successors 1803 
    -- members (2) 
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi11x_xloopexit_xx_x_crit_edgex_xix_xix_xi11_PhiReq/phi_stmt_2902/phi_stmt_2902_sources/type_cast_2908/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi11x_xloopexit_xx_x_crit_edgex_xix_xix_xi11_PhiReq/phi_stmt_2902/phi_stmt_2902_sources/type_cast_2908/SplitProtocol/Sample/ra
      -- 
    ra_17622_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2908_inst_ack_0, ack => cp_elements(1800)); -- 
    -- CP-element group 1801 transition  output  bypass 
    -- predecessors 1798 
    -- successors 1802 
    -- members (2) 
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi11x_xloopexit_xx_x_crit_edgex_xix_xix_xi11_PhiReq/phi_stmt_2902/phi_stmt_2902_sources/type_cast_2908/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi11x_xloopexit_xx_x_crit_edgex_xix_xix_xi11_PhiReq/phi_stmt_2902/phi_stmt_2902_sources/type_cast_2908/SplitProtocol/Update/cr
      -- 
    cp_elements(1801) <= cp_elements(1798);
    cr_17626_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1801), ack => type_cast_2908_inst_req_1); -- 
    -- CP-element group 1802 transition  input  bypass 
    -- predecessors 1801 
    -- successors 1803 
    -- members (2) 
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi11x_xloopexit_xx_x_crit_edgex_xix_xix_xi11_PhiReq/phi_stmt_2902/phi_stmt_2902_sources/type_cast_2908/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi11x_xloopexit_xx_x_crit_edgex_xix_xix_xi11_PhiReq/phi_stmt_2902/phi_stmt_2902_sources/type_cast_2908/SplitProtocol/Update/ca
      -- 
    ca_17627_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2908_inst_ack_1, ack => cp_elements(1802)); -- 
    -- CP-element group 1803 join  transition  output  bypass 
    -- predecessors 1800 1802 
    -- successors 1804 
    -- members (5) 
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi11x_xloopexit_xx_x_crit_edgex_xix_xix_xi11_PhiReq/phi_stmt_2902/$exit
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi11x_xloopexit_xx_x_crit_edgex_xix_xix_xi11_PhiReq/phi_stmt_2902/phi_stmt_2902_sources/$exit
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi11x_xloopexit_xx_x_crit_edgex_xix_xix_xi11_PhiReq/phi_stmt_2902/phi_stmt_2902_sources/type_cast_2908/$exit
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi11x_xloopexit_xx_x_crit_edgex_xix_xix_xi11_PhiReq/phi_stmt_2902/phi_stmt_2902_sources/type_cast_2908/SplitProtocol/$exit
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi11x_xloopexit_xx_x_crit_edgex_xix_xix_xi11_PhiReq/phi_stmt_2902/phi_stmt_2902_req
      -- 
    cp_element_group_1803: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1803"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1800) & cp_elements(1802);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1803), clk => clk, reset => reset); --
    end block;
    phi_stmt_2902_req_17628_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1803), ack => phi_stmt_2902_req_1); -- 
    -- CP-element group 1804 join  transition  bypass 
    -- predecessors 1797 1803 
    -- successors 1805 
    -- members (1) 
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi11x_xloopexit_xx_x_crit_edgex_xix_xix_xi11_PhiReq/$exit
      -- 
    cp_element_group_1804: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1804"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1797) & cp_elements(1803);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1804), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1805 merge  place  bypass 
    -- predecessors 1784 1804 
    -- successors 1806 
    -- members (1) 
      -- 	branch_block_stmt_2042/merge_stmt_2895_PhiReqMerge
      -- 
    cp_elements(1805) <= OrReduce(cp_elements(1784) & cp_elements(1804));
    -- CP-element group 1806 fork  transition  bypass 
    -- predecessors 1805 
    -- successors 1807 1808 
    -- members (1) 
      -- 	branch_block_stmt_2042/merge_stmt_2895_PhiAck/$entry
      -- 
    cp_elements(1806) <= cp_elements(1805);
    -- CP-element group 1807 transition  input  bypass 
    -- predecessors 1806 
    -- successors 1809 
    -- members (1) 
      -- 	branch_block_stmt_2042/merge_stmt_2895_PhiAck/phi_stmt_2896_ack
      -- 
    phi_stmt_2896_ack_17633_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2896_ack_0, ack => cp_elements(1807)); -- 
    -- CP-element group 1808 transition  input  bypass 
    -- predecessors 1806 
    -- successors 1809 
    -- members (1) 
      -- 	branch_block_stmt_2042/merge_stmt_2895_PhiAck/phi_stmt_2902_ack
      -- 
    phi_stmt_2902_ack_17634_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2902_ack_0, ack => cp_elements(1808)); -- 
    -- CP-element group 1809 join  transition  bypass 
    -- predecessors 1807 1808 
    -- successors 35 
    -- members (1) 
      -- 	branch_block_stmt_2042/merge_stmt_2895_PhiAck/$exit
      -- 
    cp_element_group_1809: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1809"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1807) & cp_elements(1808);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1809), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1810 transition  output  bypass 
    -- predecessors 622 
    -- successors 1811 
    -- members (2) 
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi11_xx_xloopexitx_xix_xix_xi13x_xloopexit_PhiReq/phi_stmt_2932/phi_stmt_2932_sources/type_cast_2935/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi11_xx_xloopexitx_xix_xix_xi13x_xloopexit_PhiReq/phi_stmt_2932/phi_stmt_2932_sources/type_cast_2935/SplitProtocol/Sample/rr
      -- 
    cp_elements(1810) <= cp_elements(622);
    rr_17657_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1810), ack => type_cast_2935_inst_req_0); -- 
    -- CP-element group 1811 transition  input  bypass 
    -- predecessors 1810 
    -- successors 1814 
    -- members (2) 
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi11_xx_xloopexitx_xix_xix_xi13x_xloopexit_PhiReq/phi_stmt_2932/phi_stmt_2932_sources/type_cast_2935/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi11_xx_xloopexitx_xix_xix_xi13x_xloopexit_PhiReq/phi_stmt_2932/phi_stmt_2932_sources/type_cast_2935/SplitProtocol/Sample/ra
      -- 
    ra_17658_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2935_inst_ack_0, ack => cp_elements(1811)); -- 
    -- CP-element group 1812 transition  output  bypass 
    -- predecessors 622 
    -- successors 1813 
    -- members (2) 
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi11_xx_xloopexitx_xix_xix_xi13x_xloopexit_PhiReq/phi_stmt_2932/phi_stmt_2932_sources/type_cast_2935/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi11_xx_xloopexitx_xix_xix_xi13x_xloopexit_PhiReq/phi_stmt_2932/phi_stmt_2932_sources/type_cast_2935/SplitProtocol/Update/cr
      -- 
    cp_elements(1812) <= cp_elements(622);
    cr_17662_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1812), ack => type_cast_2935_inst_req_1); -- 
    -- CP-element group 1813 transition  input  bypass 
    -- predecessors 1812 
    -- successors 1814 
    -- members (2) 
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi11_xx_xloopexitx_xix_xix_xi13x_xloopexit_PhiReq/phi_stmt_2932/phi_stmt_2932_sources/type_cast_2935/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi11_xx_xloopexitx_xix_xix_xi13x_xloopexit_PhiReq/phi_stmt_2932/phi_stmt_2932_sources/type_cast_2935/SplitProtocol/Update/ca
      -- 
    ca_17663_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2935_inst_ack_1, ack => cp_elements(1813)); -- 
    -- CP-element group 1814 join  transition  place  output  bypass 
    -- predecessors 1811 1813 
    -- successors 1815 
    -- members (8) 
      -- 	branch_block_stmt_2042/merge_stmt_2931_PhiReqMerge
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi11_xx_xloopexitx_xix_xix_xi13x_xloopexit_PhiReq/$exit
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi11_xx_xloopexitx_xix_xix_xi13x_xloopexit_PhiReq/phi_stmt_2932/$exit
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi11_xx_xloopexitx_xix_xix_xi13x_xloopexit_PhiReq/phi_stmt_2932/phi_stmt_2932_sources/$exit
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi11_xx_xloopexitx_xix_xix_xi13x_xloopexit_PhiReq/phi_stmt_2932/phi_stmt_2932_sources/type_cast_2935/$exit
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi11_xx_xloopexitx_xix_xix_xi13x_xloopexit_PhiReq/phi_stmt_2932/phi_stmt_2932_sources/type_cast_2935/SplitProtocol/$exit
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi11_xx_xloopexitx_xix_xix_xi13x_xloopexit_PhiReq/phi_stmt_2932/phi_stmt_2932_req
      -- 	branch_block_stmt_2042/merge_stmt_2931_PhiAck/$entry
      -- 
    cp_element_group_1814: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1814"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1811) & cp_elements(1813);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1814), clk => clk, reset => reset); --
    end block;
    phi_stmt_2932_req_17664_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1814), ack => phi_stmt_2932_req_0); -- 
    -- CP-element group 1815 transition  input  bypass 
    -- predecessors 1814 
    -- successors 37 
    -- members (2) 
      -- 	branch_block_stmt_2042/merge_stmt_2931_PhiAck/$exit
      -- 	branch_block_stmt_2042/merge_stmt_2931_PhiAck/phi_stmt_2932_ack
      -- 
    phi_stmt_2932_ack_17669_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2932_ack_0, ack => cp_elements(1815)); -- 
    -- CP-element group 1816 transition  bypass 
    -- predecessors 555 
    -- successors 1818 
    -- members (4) 
      -- 	branch_block_stmt_2042/bb_26_xx_xloopexitx_xix_xix_xi13_PhiReq/phi_stmt_2939/phi_stmt_2939_sources/type_cast_2945/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_2042/bb_26_xx_xloopexitx_xix_xix_xi13_PhiReq/phi_stmt_2939/phi_stmt_2939_sources/type_cast_2945/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_2042/bb_26_xx_xloopexitx_xix_xix_xi13_PhiReq/phi_stmt_2939/phi_stmt_2939_sources/type_cast_2945/SplitProtocol/Sample/rr
      -- 	branch_block_stmt_2042/bb_26_xx_xloopexitx_xix_xix_xi13_PhiReq/phi_stmt_2939/phi_stmt_2939_sources/type_cast_2945/SplitProtocol/Sample/ra
      -- 
    cp_elements(1816) <= cp_elements(555);
    -- CP-element group 1817 transition  bypass 
    -- predecessors 555 
    -- successors 1818 
    -- members (4) 
      -- 	branch_block_stmt_2042/bb_26_xx_xloopexitx_xix_xix_xi13_PhiReq/phi_stmt_2939/phi_stmt_2939_sources/type_cast_2945/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_2042/bb_26_xx_xloopexitx_xix_xix_xi13_PhiReq/phi_stmt_2939/phi_stmt_2939_sources/type_cast_2945/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_2042/bb_26_xx_xloopexitx_xix_xix_xi13_PhiReq/phi_stmt_2939/phi_stmt_2939_sources/type_cast_2945/SplitProtocol/Update/cr
      -- 	branch_block_stmt_2042/bb_26_xx_xloopexitx_xix_xix_xi13_PhiReq/phi_stmt_2939/phi_stmt_2939_sources/type_cast_2945/SplitProtocol/Update/ca
      -- 
    cp_elements(1817) <= cp_elements(555);
    -- CP-element group 1818 join  transition  output  bypass 
    -- predecessors 1816 1817 
    -- successors 1824 
    -- members (6) 
      -- 	branch_block_stmt_2042/bb_26_xx_xloopexitx_xix_xix_xi13_PhiReq/$exit
      -- 	branch_block_stmt_2042/bb_26_xx_xloopexitx_xix_xix_xi13_PhiReq/phi_stmt_2939/$exit
      -- 	branch_block_stmt_2042/bb_26_xx_xloopexitx_xix_xix_xi13_PhiReq/phi_stmt_2939/phi_stmt_2939_sources/$exit
      -- 	branch_block_stmt_2042/bb_26_xx_xloopexitx_xix_xix_xi13_PhiReq/phi_stmt_2939/phi_stmt_2939_sources/type_cast_2945/$exit
      -- 	branch_block_stmt_2042/bb_26_xx_xloopexitx_xix_xix_xi13_PhiReq/phi_stmt_2939/phi_stmt_2939_sources/type_cast_2945/SplitProtocol/$exit
      -- 	branch_block_stmt_2042/bb_26_xx_xloopexitx_xix_xix_xi13_PhiReq/phi_stmt_2939/phi_stmt_2939_req
      -- 
    cp_element_group_1818: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1818"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1816) & cp_elements(1817);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1818), clk => clk, reset => reset); --
    end block;
    phi_stmt_2939_req_17695_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1818), ack => phi_stmt_2939_req_0); -- 
    -- CP-element group 1819 transition  output  bypass 
    -- predecessors 37 
    -- successors 1820 
    -- members (2) 
      -- 	branch_block_stmt_2042/xx_xloopexitx_xix_xix_xi13x_xloopexit_xx_xloopexitx_xix_xix_xi13_PhiReq/phi_stmt_2939/phi_stmt_2939_sources/type_cast_2945/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_2042/xx_xloopexitx_xix_xix_xi13x_xloopexit_xx_xloopexitx_xix_xix_xi13_PhiReq/phi_stmt_2939/phi_stmt_2939_sources/type_cast_2945/SplitProtocol/Sample/rr
      -- 
    cp_elements(1819) <= cp_elements(37);
    rr_17714_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1819), ack => type_cast_2945_inst_req_0); -- 
    -- CP-element group 1820 transition  input  bypass 
    -- predecessors 1819 
    -- successors 1823 
    -- members (2) 
      -- 	branch_block_stmt_2042/xx_xloopexitx_xix_xix_xi13x_xloopexit_xx_xloopexitx_xix_xix_xi13_PhiReq/phi_stmt_2939/phi_stmt_2939_sources/type_cast_2945/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_2042/xx_xloopexitx_xix_xix_xi13x_xloopexit_xx_xloopexitx_xix_xix_xi13_PhiReq/phi_stmt_2939/phi_stmt_2939_sources/type_cast_2945/SplitProtocol/Sample/ra
      -- 
    ra_17715_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2945_inst_ack_0, ack => cp_elements(1820)); -- 
    -- CP-element group 1821 transition  output  bypass 
    -- predecessors 37 
    -- successors 1822 
    -- members (2) 
      -- 	branch_block_stmt_2042/xx_xloopexitx_xix_xix_xi13x_xloopexit_xx_xloopexitx_xix_xix_xi13_PhiReq/phi_stmt_2939/phi_stmt_2939_sources/type_cast_2945/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_2042/xx_xloopexitx_xix_xix_xi13x_xloopexit_xx_xloopexitx_xix_xix_xi13_PhiReq/phi_stmt_2939/phi_stmt_2939_sources/type_cast_2945/SplitProtocol/Update/cr
      -- 
    cp_elements(1821) <= cp_elements(37);
    cr_17719_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1821), ack => type_cast_2945_inst_req_1); -- 
    -- CP-element group 1822 transition  input  bypass 
    -- predecessors 1821 
    -- successors 1823 
    -- members (2) 
      -- 	branch_block_stmt_2042/xx_xloopexitx_xix_xix_xi13x_xloopexit_xx_xloopexitx_xix_xix_xi13_PhiReq/phi_stmt_2939/phi_stmt_2939_sources/type_cast_2945/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_2042/xx_xloopexitx_xix_xix_xi13x_xloopexit_xx_xloopexitx_xix_xix_xi13_PhiReq/phi_stmt_2939/phi_stmt_2939_sources/type_cast_2945/SplitProtocol/Update/ca
      -- 
    ca_17720_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2945_inst_ack_1, ack => cp_elements(1822)); -- 
    -- CP-element group 1823 join  transition  output  bypass 
    -- predecessors 1820 1822 
    -- successors 1824 
    -- members (6) 
      -- 	branch_block_stmt_2042/xx_xloopexitx_xix_xix_xi13x_xloopexit_xx_xloopexitx_xix_xix_xi13_PhiReq/$exit
      -- 	branch_block_stmt_2042/xx_xloopexitx_xix_xix_xi13x_xloopexit_xx_xloopexitx_xix_xix_xi13_PhiReq/phi_stmt_2939/$exit
      -- 	branch_block_stmt_2042/xx_xloopexitx_xix_xix_xi13x_xloopexit_xx_xloopexitx_xix_xix_xi13_PhiReq/phi_stmt_2939/phi_stmt_2939_sources/$exit
      -- 	branch_block_stmt_2042/xx_xloopexitx_xix_xix_xi13x_xloopexit_xx_xloopexitx_xix_xix_xi13_PhiReq/phi_stmt_2939/phi_stmt_2939_sources/type_cast_2945/$exit
      -- 	branch_block_stmt_2042/xx_xloopexitx_xix_xix_xi13x_xloopexit_xx_xloopexitx_xix_xix_xi13_PhiReq/phi_stmt_2939/phi_stmt_2939_sources/type_cast_2945/SplitProtocol/$exit
      -- 	branch_block_stmt_2042/xx_xloopexitx_xix_xix_xi13x_xloopexit_xx_xloopexitx_xix_xix_xi13_PhiReq/phi_stmt_2939/phi_stmt_2939_req
      -- 
    cp_element_group_1823: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1823"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1820) & cp_elements(1822);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1823), clk => clk, reset => reset); --
    end block;
    phi_stmt_2939_req_17721_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1823), ack => phi_stmt_2939_req_1); -- 
    -- CP-element group 1824 merge  place  bypass 
    -- predecessors 1818 1823 
    -- successors 1825 
    -- members (1) 
      -- 	branch_block_stmt_2042/merge_stmt_2938_PhiReqMerge
      -- 
    cp_elements(1824) <= OrReduce(cp_elements(1818) & cp_elements(1823));
    -- CP-element group 1825 transition  bypass 
    -- predecessors 1824 
    -- successors 1826 
    -- members (1) 
      -- 	branch_block_stmt_2042/merge_stmt_2938_PhiAck/$entry
      -- 
    cp_elements(1825) <= cp_elements(1824);
    -- CP-element group 1826 fork  transition  place  input  bypass 
    -- predecessors 1825 
    -- successors 1838 1844 
    -- members (7) 
      -- 	branch_block_stmt_2042/xx_xloopexitx_xix_xix_xi13_udiv32x_xexitx_xpreheaderx_xix_xi16
      -- 	branch_block_stmt_2042/merge_stmt_2938__exit__
      -- 	branch_block_stmt_2042/merge_stmt_2938_PhiAck/$exit
      -- 	branch_block_stmt_2042/merge_stmt_2938_PhiAck/phi_stmt_2939_ack
      -- 	branch_block_stmt_2042/xx_xloopexitx_xix_xix_xi13_udiv32x_xexitx_xpreheaderx_xix_xi16_PhiReq/$entry
      -- 	branch_block_stmt_2042/xx_xloopexitx_xix_xix_xi13_udiv32x_xexitx_xpreheaderx_xix_xi16_PhiReq/phi_stmt_2949/$entry
      -- 	branch_block_stmt_2042/xx_xloopexitx_xix_xix_xi13_udiv32x_xexitx_xpreheaderx_xix_xi16_PhiReq/phi_stmt_2949/phi_stmt_2949_sources/$entry
      -- 
    phi_stmt_2939_ack_17726_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2939_ack_0, ack => cp_elements(1826)); -- 
    -- CP-element group 1827 fork  transition  bypass 
    -- predecessors 557 
    -- successors 1828 1829 
    -- members (2) 
      -- 	branch_block_stmt_2042/bb_26_udiv32x_xexitx_xpreheaderx_xix_xi16_PhiReq/phi_stmt_2949/phi_stmt_2949_sources/type_cast_2952/$entry
      -- 	branch_block_stmt_2042/bb_26_udiv32x_xexitx_xpreheaderx_xix_xi16_PhiReq/phi_stmt_2949/phi_stmt_2949_sources/type_cast_2952/SplitProtocol/$entry
      -- 
    cp_elements(1827) <= cp_elements(557);
    -- CP-element group 1828 transition  bypass 
    -- predecessors 1827 
    -- successors 1830 
    -- members (4) 
      -- 	branch_block_stmt_2042/bb_26_udiv32x_xexitx_xpreheaderx_xix_xi16_PhiReq/phi_stmt_2949/phi_stmt_2949_sources/type_cast_2952/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_2042/bb_26_udiv32x_xexitx_xpreheaderx_xix_xi16_PhiReq/phi_stmt_2949/phi_stmt_2949_sources/type_cast_2952/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_2042/bb_26_udiv32x_xexitx_xpreheaderx_xix_xi16_PhiReq/phi_stmt_2949/phi_stmt_2949_sources/type_cast_2952/SplitProtocol/Sample/rr
      -- 	branch_block_stmt_2042/bb_26_udiv32x_xexitx_xpreheaderx_xix_xi16_PhiReq/phi_stmt_2949/phi_stmt_2949_sources/type_cast_2952/SplitProtocol/Sample/ra
      -- 
    cp_elements(1828) <= cp_elements(1827);
    -- CP-element group 1829 transition  bypass 
    -- predecessors 1827 
    -- successors 1830 
    -- members (4) 
      -- 	branch_block_stmt_2042/bb_26_udiv32x_xexitx_xpreheaderx_xix_xi16_PhiReq/phi_stmt_2949/phi_stmt_2949_sources/type_cast_2952/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_2042/bb_26_udiv32x_xexitx_xpreheaderx_xix_xi16_PhiReq/phi_stmt_2949/phi_stmt_2949_sources/type_cast_2952/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_2042/bb_26_udiv32x_xexitx_xpreheaderx_xix_xi16_PhiReq/phi_stmt_2949/phi_stmt_2949_sources/type_cast_2952/SplitProtocol/Update/cr
      -- 	branch_block_stmt_2042/bb_26_udiv32x_xexitx_xpreheaderx_xix_xi16_PhiReq/phi_stmt_2949/phi_stmt_2949_sources/type_cast_2952/SplitProtocol/Update/ca
      -- 
    cp_elements(1829) <= cp_elements(1827);
    -- CP-element group 1830 join  transition  bypass 
    -- predecessors 1828 1829 
    -- successors 1837 
    -- members (2) 
      -- 	branch_block_stmt_2042/bb_26_udiv32x_xexitx_xpreheaderx_xix_xi16_PhiReq/phi_stmt_2949/phi_stmt_2949_sources/type_cast_2952/$exit
      -- 	branch_block_stmt_2042/bb_26_udiv32x_xexitx_xpreheaderx_xix_xi16_PhiReq/phi_stmt_2949/phi_stmt_2949_sources/type_cast_2952/SplitProtocol/$exit
      -- 
    cp_element_group_1830: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1830"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1828) & cp_elements(1829);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1830), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1831 fork  transition  bypass 
    -- predecessors 557 
    -- successors 1832 1834 
    -- members (2) 
      -- 	branch_block_stmt_2042/bb_26_udiv32x_xexitx_xpreheaderx_xix_xi16_PhiReq/phi_stmt_2949/phi_stmt_2949_sources/type_cast_2954/$entry
      -- 	branch_block_stmt_2042/bb_26_udiv32x_xexitx_xpreheaderx_xix_xi16_PhiReq/phi_stmt_2949/phi_stmt_2949_sources/type_cast_2954/SplitProtocol/$entry
      -- 
    cp_elements(1831) <= cp_elements(557);
    -- CP-element group 1832 transition  output  bypass 
    -- predecessors 1831 
    -- successors 1833 
    -- members (2) 
      -- 	branch_block_stmt_2042/bb_26_udiv32x_xexitx_xpreheaderx_xix_xi16_PhiReq/phi_stmt_2949/phi_stmt_2949_sources/type_cast_2954/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_2042/bb_26_udiv32x_xexitx_xpreheaderx_xix_xi16_PhiReq/phi_stmt_2949/phi_stmt_2949_sources/type_cast_2954/SplitProtocol/Sample/rr
      -- 
    cp_elements(1832) <= cp_elements(1831);
    rr_17761_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1832), ack => type_cast_2954_inst_req_0); -- 
    -- CP-element group 1833 transition  input  bypass 
    -- predecessors 1832 
    -- successors 1836 
    -- members (2) 
      -- 	branch_block_stmt_2042/bb_26_udiv32x_xexitx_xpreheaderx_xix_xi16_PhiReq/phi_stmt_2949/phi_stmt_2949_sources/type_cast_2954/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_2042/bb_26_udiv32x_xexitx_xpreheaderx_xix_xi16_PhiReq/phi_stmt_2949/phi_stmt_2949_sources/type_cast_2954/SplitProtocol/Sample/ra
      -- 
    ra_17762_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2954_inst_ack_0, ack => cp_elements(1833)); -- 
    -- CP-element group 1834 transition  output  bypass 
    -- predecessors 1831 
    -- successors 1835 
    -- members (2) 
      -- 	branch_block_stmt_2042/bb_26_udiv32x_xexitx_xpreheaderx_xix_xi16_PhiReq/phi_stmt_2949/phi_stmt_2949_sources/type_cast_2954/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_2042/bb_26_udiv32x_xexitx_xpreheaderx_xix_xi16_PhiReq/phi_stmt_2949/phi_stmt_2949_sources/type_cast_2954/SplitProtocol/Update/cr
      -- 
    cp_elements(1834) <= cp_elements(1831);
    cr_17766_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1834), ack => type_cast_2954_inst_req_1); -- 
    -- CP-element group 1835 transition  input  bypass 
    -- predecessors 1834 
    -- successors 1836 
    -- members (2) 
      -- 	branch_block_stmt_2042/bb_26_udiv32x_xexitx_xpreheaderx_xix_xi16_PhiReq/phi_stmt_2949/phi_stmt_2949_sources/type_cast_2954/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_2042/bb_26_udiv32x_xexitx_xpreheaderx_xix_xi16_PhiReq/phi_stmt_2949/phi_stmt_2949_sources/type_cast_2954/SplitProtocol/Update/ca
      -- 
    ca_17767_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2954_inst_ack_1, ack => cp_elements(1835)); -- 
    -- CP-element group 1836 join  transition  bypass 
    -- predecessors 1833 1835 
    -- successors 1837 
    -- members (2) 
      -- 	branch_block_stmt_2042/bb_26_udiv32x_xexitx_xpreheaderx_xix_xi16_PhiReq/phi_stmt_2949/phi_stmt_2949_sources/type_cast_2954/$exit
      -- 	branch_block_stmt_2042/bb_26_udiv32x_xexitx_xpreheaderx_xix_xi16_PhiReq/phi_stmt_2949/phi_stmt_2949_sources/type_cast_2954/SplitProtocol/$exit
      -- 
    cp_element_group_1836: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1836"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1833) & cp_elements(1835);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1836), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1837 join  transition  output  bypass 
    -- predecessors 1830 1836 
    -- successors 1849 
    -- members (4) 
      -- 	branch_block_stmt_2042/bb_26_udiv32x_xexitx_xpreheaderx_xix_xi16_PhiReq/$exit
      -- 	branch_block_stmt_2042/bb_26_udiv32x_xexitx_xpreheaderx_xix_xi16_PhiReq/phi_stmt_2949/$exit
      -- 	branch_block_stmt_2042/bb_26_udiv32x_xexitx_xpreheaderx_xix_xi16_PhiReq/phi_stmt_2949/phi_stmt_2949_sources/$exit
      -- 	branch_block_stmt_2042/bb_26_udiv32x_xexitx_xpreheaderx_xix_xi16_PhiReq/phi_stmt_2949/phi_stmt_2949_req
      -- 
    cp_element_group_1837: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1837"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1830) & cp_elements(1836);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1837), clk => clk, reset => reset); --
    end block;
    phi_stmt_2949_req_17768_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1837), ack => phi_stmt_2949_req_1); -- 
    -- CP-element group 1838 fork  transition  bypass 
    -- predecessors 1826 
    -- successors 1839 1841 
    -- members (2) 
      -- 	branch_block_stmt_2042/xx_xloopexitx_xix_xix_xi13_udiv32x_xexitx_xpreheaderx_xix_xi16_PhiReq/phi_stmt_2949/phi_stmt_2949_sources/type_cast_2952/$entry
      -- 	branch_block_stmt_2042/xx_xloopexitx_xix_xix_xi13_udiv32x_xexitx_xpreheaderx_xix_xi16_PhiReq/phi_stmt_2949/phi_stmt_2949_sources/type_cast_2952/SplitProtocol/$entry
      -- 
    cp_elements(1838) <= cp_elements(1826);
    -- CP-element group 1839 transition  output  bypass 
    -- predecessors 1838 
    -- successors 1840 
    -- members (2) 
      -- 	branch_block_stmt_2042/xx_xloopexitx_xix_xix_xi13_udiv32x_xexitx_xpreheaderx_xix_xi16_PhiReq/phi_stmt_2949/phi_stmt_2949_sources/type_cast_2952/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_2042/xx_xloopexitx_xix_xix_xi13_udiv32x_xexitx_xpreheaderx_xix_xi16_PhiReq/phi_stmt_2949/phi_stmt_2949_sources/type_cast_2952/SplitProtocol/Sample/rr
      -- 
    cp_elements(1839) <= cp_elements(1838);
    rr_17787_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1839), ack => type_cast_2952_inst_req_0); -- 
    -- CP-element group 1840 transition  input  bypass 
    -- predecessors 1839 
    -- successors 1843 
    -- members (2) 
      -- 	branch_block_stmt_2042/xx_xloopexitx_xix_xix_xi13_udiv32x_xexitx_xpreheaderx_xix_xi16_PhiReq/phi_stmt_2949/phi_stmt_2949_sources/type_cast_2952/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_2042/xx_xloopexitx_xix_xix_xi13_udiv32x_xexitx_xpreheaderx_xix_xi16_PhiReq/phi_stmt_2949/phi_stmt_2949_sources/type_cast_2952/SplitProtocol/Sample/ra
      -- 
    ra_17788_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2952_inst_ack_0, ack => cp_elements(1840)); -- 
    -- CP-element group 1841 transition  output  bypass 
    -- predecessors 1838 
    -- successors 1842 
    -- members (2) 
      -- 	branch_block_stmt_2042/xx_xloopexitx_xix_xix_xi13_udiv32x_xexitx_xpreheaderx_xix_xi16_PhiReq/phi_stmt_2949/phi_stmt_2949_sources/type_cast_2952/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_2042/xx_xloopexitx_xix_xix_xi13_udiv32x_xexitx_xpreheaderx_xix_xi16_PhiReq/phi_stmt_2949/phi_stmt_2949_sources/type_cast_2952/SplitProtocol/Update/cr
      -- 
    cp_elements(1841) <= cp_elements(1838);
    cr_17792_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1841), ack => type_cast_2952_inst_req_1); -- 
    -- CP-element group 1842 transition  input  bypass 
    -- predecessors 1841 
    -- successors 1843 
    -- members (2) 
      -- 	branch_block_stmt_2042/xx_xloopexitx_xix_xix_xi13_udiv32x_xexitx_xpreheaderx_xix_xi16_PhiReq/phi_stmt_2949/phi_stmt_2949_sources/type_cast_2952/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_2042/xx_xloopexitx_xix_xix_xi13_udiv32x_xexitx_xpreheaderx_xix_xi16_PhiReq/phi_stmt_2949/phi_stmt_2949_sources/type_cast_2952/SplitProtocol/Update/ca
      -- 
    ca_17793_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2952_inst_ack_1, ack => cp_elements(1842)); -- 
    -- CP-element group 1843 join  transition  bypass 
    -- predecessors 1840 1842 
    -- successors 1848 
    -- members (2) 
      -- 	branch_block_stmt_2042/xx_xloopexitx_xix_xix_xi13_udiv32x_xexitx_xpreheaderx_xix_xi16_PhiReq/phi_stmt_2949/phi_stmt_2949_sources/type_cast_2952/$exit
      -- 	branch_block_stmt_2042/xx_xloopexitx_xix_xix_xi13_udiv32x_xexitx_xpreheaderx_xix_xi16_PhiReq/phi_stmt_2949/phi_stmt_2949_sources/type_cast_2952/SplitProtocol/$exit
      -- 
    cp_element_group_1843: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1843"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1840) & cp_elements(1842);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1843), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1844 fork  transition  bypass 
    -- predecessors 1826 
    -- successors 1845 1846 
    -- members (2) 
      -- 	branch_block_stmt_2042/xx_xloopexitx_xix_xix_xi13_udiv32x_xexitx_xpreheaderx_xix_xi16_PhiReq/phi_stmt_2949/phi_stmt_2949_sources/type_cast_2954/$entry
      -- 	branch_block_stmt_2042/xx_xloopexitx_xix_xix_xi13_udiv32x_xexitx_xpreheaderx_xix_xi16_PhiReq/phi_stmt_2949/phi_stmt_2949_sources/type_cast_2954/SplitProtocol/$entry
      -- 
    cp_elements(1844) <= cp_elements(1826);
    -- CP-element group 1845 transition  bypass 
    -- predecessors 1844 
    -- successors 1847 
    -- members (4) 
      -- 	branch_block_stmt_2042/xx_xloopexitx_xix_xix_xi13_udiv32x_xexitx_xpreheaderx_xix_xi16_PhiReq/phi_stmt_2949/phi_stmt_2949_sources/type_cast_2954/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_2042/xx_xloopexitx_xix_xix_xi13_udiv32x_xexitx_xpreheaderx_xix_xi16_PhiReq/phi_stmt_2949/phi_stmt_2949_sources/type_cast_2954/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_2042/xx_xloopexitx_xix_xix_xi13_udiv32x_xexitx_xpreheaderx_xix_xi16_PhiReq/phi_stmt_2949/phi_stmt_2949_sources/type_cast_2954/SplitProtocol/Sample/rr
      -- 	branch_block_stmt_2042/xx_xloopexitx_xix_xix_xi13_udiv32x_xexitx_xpreheaderx_xix_xi16_PhiReq/phi_stmt_2949/phi_stmt_2949_sources/type_cast_2954/SplitProtocol/Sample/ra
      -- 
    cp_elements(1845) <= cp_elements(1844);
    -- CP-element group 1846 transition  bypass 
    -- predecessors 1844 
    -- successors 1847 
    -- members (4) 
      -- 	branch_block_stmt_2042/xx_xloopexitx_xix_xix_xi13_udiv32x_xexitx_xpreheaderx_xix_xi16_PhiReq/phi_stmt_2949/phi_stmt_2949_sources/type_cast_2954/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_2042/xx_xloopexitx_xix_xix_xi13_udiv32x_xexitx_xpreheaderx_xix_xi16_PhiReq/phi_stmt_2949/phi_stmt_2949_sources/type_cast_2954/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_2042/xx_xloopexitx_xix_xix_xi13_udiv32x_xexitx_xpreheaderx_xix_xi16_PhiReq/phi_stmt_2949/phi_stmt_2949_sources/type_cast_2954/SplitProtocol/Update/cr
      -- 	branch_block_stmt_2042/xx_xloopexitx_xix_xix_xi13_udiv32x_xexitx_xpreheaderx_xix_xi16_PhiReq/phi_stmt_2949/phi_stmt_2949_sources/type_cast_2954/SplitProtocol/Update/ca
      -- 
    cp_elements(1846) <= cp_elements(1844);
    -- CP-element group 1847 join  transition  bypass 
    -- predecessors 1845 1846 
    -- successors 1848 
    -- members (2) 
      -- 	branch_block_stmt_2042/xx_xloopexitx_xix_xix_xi13_udiv32x_xexitx_xpreheaderx_xix_xi16_PhiReq/phi_stmt_2949/phi_stmt_2949_sources/type_cast_2954/$exit
      -- 	branch_block_stmt_2042/xx_xloopexitx_xix_xix_xi13_udiv32x_xexitx_xpreheaderx_xix_xi16_PhiReq/phi_stmt_2949/phi_stmt_2949_sources/type_cast_2954/SplitProtocol/$exit
      -- 
    cp_element_group_1847: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1847"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1845) & cp_elements(1846);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1847), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1848 join  transition  output  bypass 
    -- predecessors 1843 1847 
    -- successors 1849 
    -- members (4) 
      -- 	branch_block_stmt_2042/xx_xloopexitx_xix_xix_xi13_udiv32x_xexitx_xpreheaderx_xix_xi16_PhiReq/$exit
      -- 	branch_block_stmt_2042/xx_xloopexitx_xix_xix_xi13_udiv32x_xexitx_xpreheaderx_xix_xi16_PhiReq/phi_stmt_2949/$exit
      -- 	branch_block_stmt_2042/xx_xloopexitx_xix_xix_xi13_udiv32x_xexitx_xpreheaderx_xix_xi16_PhiReq/phi_stmt_2949/phi_stmt_2949_sources/$exit
      -- 	branch_block_stmt_2042/xx_xloopexitx_xix_xix_xi13_udiv32x_xexitx_xpreheaderx_xix_xi16_PhiReq/phi_stmt_2949/phi_stmt_2949_req
      -- 
    cp_element_group_1848: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1848"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1843) & cp_elements(1847);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1848), clk => clk, reset => reset); --
    end block;
    phi_stmt_2949_req_17810_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1848), ack => phi_stmt_2949_req_0); -- 
    -- CP-element group 1849 merge  place  bypass 
    -- predecessors 1837 1848 
    -- successors 1850 
    -- members (1) 
      -- 	branch_block_stmt_2042/merge_stmt_2948_PhiReqMerge
      -- 
    cp_elements(1849) <= OrReduce(cp_elements(1837) & cp_elements(1848));
    -- CP-element group 1850 transition  bypass 
    -- predecessors 1849 
    -- successors 1851 
    -- members (1) 
      -- 	branch_block_stmt_2042/merge_stmt_2948_PhiAck/$entry
      -- 
    cp_elements(1850) <= cp_elements(1849);
    -- CP-element group 1851 transition  place  input  bypass 
    -- predecessors 1850 
    -- successors 625 
    -- members (4) 
      -- 	branch_block_stmt_2042/assign_stmt_2961_to_assign_stmt_2980__entry__
      -- 	branch_block_stmt_2042/merge_stmt_2948__exit__
      -- 	branch_block_stmt_2042/merge_stmt_2948_PhiAck/$exit
      -- 	branch_block_stmt_2042/merge_stmt_2948_PhiAck/phi_stmt_2949_ack
      -- 
    phi_stmt_2949_ack_17815_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2949_ack_0, ack => cp_elements(1851)); -- 
    -- CP-element group 1852 fork  transition  bypass 
    -- predecessors 681 
    -- successors 1853 1859 
    -- members (1) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi20_udiv32x_xexitx_xix_xi20_PhiReq/$entry
      -- 
    cp_elements(1852) <= cp_elements(681);
    -- CP-element group 1853 fork  transition  bypass 
    -- predecessors 1852 
    -- successors 1854 1856 
    -- members (4) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi20_udiv32x_xexitx_xix_xi20_PhiReq/phi_stmt_2990/$entry
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi20_udiv32x_xexitx_xix_xi20_PhiReq/phi_stmt_2990/phi_stmt_2990_sources/$entry
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi20_udiv32x_xexitx_xix_xi20_PhiReq/phi_stmt_2990/phi_stmt_2990_sources/type_cast_2993/$entry
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi20_udiv32x_xexitx_xix_xi20_PhiReq/phi_stmt_2990/phi_stmt_2990_sources/type_cast_2993/SplitProtocol/$entry
      -- 
    cp_elements(1853) <= cp_elements(1852);
    -- CP-element group 1854 transition  output  bypass 
    -- predecessors 1853 
    -- successors 1855 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi20_udiv32x_xexitx_xix_xi20_PhiReq/phi_stmt_2990/phi_stmt_2990_sources/type_cast_2993/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi20_udiv32x_xexitx_xix_xi20_PhiReq/phi_stmt_2990/phi_stmt_2990_sources/type_cast_2993/SplitProtocol/Sample/rr
      -- 
    cp_elements(1854) <= cp_elements(1853);
    rr_17846_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1854), ack => type_cast_2993_inst_req_0); -- 
    -- CP-element group 1855 transition  input  bypass 
    -- predecessors 1854 
    -- successors 1858 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi20_udiv32x_xexitx_xix_xi20_PhiReq/phi_stmt_2990/phi_stmt_2990_sources/type_cast_2993/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi20_udiv32x_xexitx_xix_xi20_PhiReq/phi_stmt_2990/phi_stmt_2990_sources/type_cast_2993/SplitProtocol/Sample/ra
      -- 
    ra_17847_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2993_inst_ack_0, ack => cp_elements(1855)); -- 
    -- CP-element group 1856 transition  output  bypass 
    -- predecessors 1853 
    -- successors 1857 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi20_udiv32x_xexitx_xix_xi20_PhiReq/phi_stmt_2990/phi_stmt_2990_sources/type_cast_2993/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi20_udiv32x_xexitx_xix_xi20_PhiReq/phi_stmt_2990/phi_stmt_2990_sources/type_cast_2993/SplitProtocol/Update/cr
      -- 
    cp_elements(1856) <= cp_elements(1853);
    cr_17851_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1856), ack => type_cast_2993_inst_req_1); -- 
    -- CP-element group 1857 transition  input  bypass 
    -- predecessors 1856 
    -- successors 1858 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi20_udiv32x_xexitx_xix_xi20_PhiReq/phi_stmt_2990/phi_stmt_2990_sources/type_cast_2993/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi20_udiv32x_xexitx_xix_xi20_PhiReq/phi_stmt_2990/phi_stmt_2990_sources/type_cast_2993/SplitProtocol/Update/ca
      -- 
    ca_17852_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2993_inst_ack_1, ack => cp_elements(1857)); -- 
    -- CP-element group 1858 join  transition  output  bypass 
    -- predecessors 1855 1857 
    -- successors 1871 
    -- members (5) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi20_udiv32x_xexitx_xix_xi20_PhiReq/phi_stmt_2990/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi20_udiv32x_xexitx_xix_xi20_PhiReq/phi_stmt_2990/phi_stmt_2990_sources/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi20_udiv32x_xexitx_xix_xi20_PhiReq/phi_stmt_2990/phi_stmt_2990_sources/type_cast_2993/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi20_udiv32x_xexitx_xix_xi20_PhiReq/phi_stmt_2990/phi_stmt_2990_sources/type_cast_2993/SplitProtocol/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi20_udiv32x_xexitx_xix_xi20_PhiReq/phi_stmt_2990/phi_stmt_2990_req
      -- 
    cp_element_group_1858: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1858"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1855) & cp_elements(1857);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1858), clk => clk, reset => reset); --
    end block;
    phi_stmt_2990_req_17853_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1858), ack => phi_stmt_2990_req_0); -- 
    -- CP-element group 1859 fork  transition  bypass 
    -- predecessors 1852 
    -- successors 1860 1866 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi20_udiv32x_xexitx_xix_xi20_PhiReq/phi_stmt_2997/$entry
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi20_udiv32x_xexitx_xix_xi20_PhiReq/phi_stmt_2997/phi_stmt_2997_sources/$entry
      -- 
    cp_elements(1859) <= cp_elements(1852);
    -- CP-element group 1860 fork  transition  bypass 
    -- predecessors 1859 
    -- successors 1861 1863 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi20_udiv32x_xexitx_xix_xi20_PhiReq/phi_stmt_2997/phi_stmt_2997_sources/type_cast_3000/$entry
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi20_udiv32x_xexitx_xix_xi20_PhiReq/phi_stmt_2997/phi_stmt_2997_sources/type_cast_3000/SplitProtocol/$entry
      -- 
    cp_elements(1860) <= cp_elements(1859);
    -- CP-element group 1861 transition  output  bypass 
    -- predecessors 1860 
    -- successors 1862 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi20_udiv32x_xexitx_xix_xi20_PhiReq/phi_stmt_2997/phi_stmt_2997_sources/type_cast_3000/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi20_udiv32x_xexitx_xix_xi20_PhiReq/phi_stmt_2997/phi_stmt_2997_sources/type_cast_3000/SplitProtocol/Sample/rr
      -- 
    cp_elements(1861) <= cp_elements(1860);
    rr_17869_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1861), ack => type_cast_3000_inst_req_0); -- 
    -- CP-element group 1862 transition  input  bypass 
    -- predecessors 1861 
    -- successors 1865 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi20_udiv32x_xexitx_xix_xi20_PhiReq/phi_stmt_2997/phi_stmt_2997_sources/type_cast_3000/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi20_udiv32x_xexitx_xix_xi20_PhiReq/phi_stmt_2997/phi_stmt_2997_sources/type_cast_3000/SplitProtocol/Sample/ra
      -- 
    ra_17870_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3000_inst_ack_0, ack => cp_elements(1862)); -- 
    -- CP-element group 1863 transition  output  bypass 
    -- predecessors 1860 
    -- successors 1864 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi20_udiv32x_xexitx_xix_xi20_PhiReq/phi_stmt_2997/phi_stmt_2997_sources/type_cast_3000/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi20_udiv32x_xexitx_xix_xi20_PhiReq/phi_stmt_2997/phi_stmt_2997_sources/type_cast_3000/SplitProtocol/Update/cr
      -- 
    cp_elements(1863) <= cp_elements(1860);
    cr_17874_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1863), ack => type_cast_3000_inst_req_1); -- 
    -- CP-element group 1864 transition  input  bypass 
    -- predecessors 1863 
    -- successors 1865 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi20_udiv32x_xexitx_xix_xi20_PhiReq/phi_stmt_2997/phi_stmt_2997_sources/type_cast_3000/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi20_udiv32x_xexitx_xix_xi20_PhiReq/phi_stmt_2997/phi_stmt_2997_sources/type_cast_3000/SplitProtocol/Update/ca
      -- 
    ca_17875_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3000_inst_ack_1, ack => cp_elements(1864)); -- 
    -- CP-element group 1865 join  transition  bypass 
    -- predecessors 1862 1864 
    -- successors 1870 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi20_udiv32x_xexitx_xix_xi20_PhiReq/phi_stmt_2997/phi_stmt_2997_sources/type_cast_3000/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi20_udiv32x_xexitx_xix_xi20_PhiReq/phi_stmt_2997/phi_stmt_2997_sources/type_cast_3000/SplitProtocol/$exit
      -- 
    cp_element_group_1865: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1865"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1862) & cp_elements(1864);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1865), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1866 fork  transition  bypass 
    -- predecessors 1859 
    -- successors 1867 1868 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi20_udiv32x_xexitx_xix_xi20_PhiReq/phi_stmt_2997/phi_stmt_2997_sources/type_cast_3002/$entry
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi20_udiv32x_xexitx_xix_xi20_PhiReq/phi_stmt_2997/phi_stmt_2997_sources/type_cast_3002/SplitProtocol/$entry
      -- 
    cp_elements(1866) <= cp_elements(1859);
    -- CP-element group 1867 transition  bypass 
    -- predecessors 1866 
    -- successors 1869 
    -- members (4) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi20_udiv32x_xexitx_xix_xi20_PhiReq/phi_stmt_2997/phi_stmt_2997_sources/type_cast_3002/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi20_udiv32x_xexitx_xix_xi20_PhiReq/phi_stmt_2997/phi_stmt_2997_sources/type_cast_3002/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi20_udiv32x_xexitx_xix_xi20_PhiReq/phi_stmt_2997/phi_stmt_2997_sources/type_cast_3002/SplitProtocol/Sample/rr
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi20_udiv32x_xexitx_xix_xi20_PhiReq/phi_stmt_2997/phi_stmt_2997_sources/type_cast_3002/SplitProtocol/Sample/ra
      -- 
    cp_elements(1867) <= cp_elements(1866);
    -- CP-element group 1868 transition  bypass 
    -- predecessors 1866 
    -- successors 1869 
    -- members (4) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi20_udiv32x_xexitx_xix_xi20_PhiReq/phi_stmt_2997/phi_stmt_2997_sources/type_cast_3002/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi20_udiv32x_xexitx_xix_xi20_PhiReq/phi_stmt_2997/phi_stmt_2997_sources/type_cast_3002/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi20_udiv32x_xexitx_xix_xi20_PhiReq/phi_stmt_2997/phi_stmt_2997_sources/type_cast_3002/SplitProtocol/Update/cr
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi20_udiv32x_xexitx_xix_xi20_PhiReq/phi_stmt_2997/phi_stmt_2997_sources/type_cast_3002/SplitProtocol/Update/ca
      -- 
    cp_elements(1868) <= cp_elements(1866);
    -- CP-element group 1869 join  transition  bypass 
    -- predecessors 1867 1868 
    -- successors 1870 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi20_udiv32x_xexitx_xix_xi20_PhiReq/phi_stmt_2997/phi_stmt_2997_sources/type_cast_3002/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi20_udiv32x_xexitx_xix_xi20_PhiReq/phi_stmt_2997/phi_stmt_2997_sources/type_cast_3002/SplitProtocol/$exit
      -- 
    cp_element_group_1869: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1869"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1867) & cp_elements(1868);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1869), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1870 join  transition  output  bypass 
    -- predecessors 1865 1869 
    -- successors 1871 
    -- members (3) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi20_udiv32x_xexitx_xix_xi20_PhiReq/phi_stmt_2997/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi20_udiv32x_xexitx_xix_xi20_PhiReq/phi_stmt_2997/phi_stmt_2997_sources/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi20_udiv32x_xexitx_xix_xi20_PhiReq/phi_stmt_2997/phi_stmt_2997_req
      -- 
    cp_element_group_1870: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1870"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1865) & cp_elements(1869);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1870), clk => clk, reset => reset); --
    end block;
    phi_stmt_2997_req_17892_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1870), ack => phi_stmt_2997_req_0); -- 
    -- CP-element group 1871 join  transition  bypass 
    -- predecessors 1858 1870 
    -- successors 1890 
    -- members (1) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi20_udiv32x_xexitx_xix_xi20_PhiReq/$exit
      -- 
    cp_element_group_1871: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1871"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1858) & cp_elements(1870);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1871), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1872 fork  transition  bypass 
    -- predecessors 38 
    -- successors 1873 1877 
    -- members (1) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi20x_xpreheader_udiv32x_xexitx_xix_xi20_PhiReq/$entry
      -- 
    cp_elements(1872) <= cp_elements(38);
    -- CP-element group 1873 fork  transition  bypass 
    -- predecessors 1872 
    -- successors 1874 1875 
    -- members (4) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi20x_xpreheader_udiv32x_xexitx_xix_xi20_PhiReq/phi_stmt_2990/$entry
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi20x_xpreheader_udiv32x_xexitx_xix_xi20_PhiReq/phi_stmt_2990/phi_stmt_2990_sources/$entry
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi20x_xpreheader_udiv32x_xexitx_xix_xi20_PhiReq/phi_stmt_2990/phi_stmt_2990_sources/type_cast_2993/$entry
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi20x_xpreheader_udiv32x_xexitx_xix_xi20_PhiReq/phi_stmt_2990/phi_stmt_2990_sources/type_cast_2993/SplitProtocol/$entry
      -- 
    cp_elements(1873) <= cp_elements(1872);
    -- CP-element group 1874 transition  bypass 
    -- predecessors 1873 
    -- successors 1876 
    -- members (4) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi20x_xpreheader_udiv32x_xexitx_xix_xi20_PhiReq/phi_stmt_2990/phi_stmt_2990_sources/type_cast_2993/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi20x_xpreheader_udiv32x_xexitx_xix_xi20_PhiReq/phi_stmt_2990/phi_stmt_2990_sources/type_cast_2993/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi20x_xpreheader_udiv32x_xexitx_xix_xi20_PhiReq/phi_stmt_2990/phi_stmt_2990_sources/type_cast_2993/SplitProtocol/Sample/rr
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi20x_xpreheader_udiv32x_xexitx_xix_xi20_PhiReq/phi_stmt_2990/phi_stmt_2990_sources/type_cast_2993/SplitProtocol/Sample/ra
      -- 
    cp_elements(1874) <= cp_elements(1873);
    -- CP-element group 1875 transition  bypass 
    -- predecessors 1873 
    -- successors 1876 
    -- members (4) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi20x_xpreheader_udiv32x_xexitx_xix_xi20_PhiReq/phi_stmt_2990/phi_stmt_2990_sources/type_cast_2993/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi20x_xpreheader_udiv32x_xexitx_xix_xi20_PhiReq/phi_stmt_2990/phi_stmt_2990_sources/type_cast_2993/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi20x_xpreheader_udiv32x_xexitx_xix_xi20_PhiReq/phi_stmt_2990/phi_stmt_2990_sources/type_cast_2993/SplitProtocol/Update/cr
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi20x_xpreheader_udiv32x_xexitx_xix_xi20_PhiReq/phi_stmt_2990/phi_stmt_2990_sources/type_cast_2993/SplitProtocol/Update/ca
      -- 
    cp_elements(1875) <= cp_elements(1873);
    -- CP-element group 1876 join  transition  output  bypass 
    -- predecessors 1874 1875 
    -- successors 1889 
    -- members (5) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi20x_xpreheader_udiv32x_xexitx_xix_xi20_PhiReq/phi_stmt_2990/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi20x_xpreheader_udiv32x_xexitx_xix_xi20_PhiReq/phi_stmt_2990/phi_stmt_2990_sources/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi20x_xpreheader_udiv32x_xexitx_xix_xi20_PhiReq/phi_stmt_2990/phi_stmt_2990_sources/type_cast_2993/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi20x_xpreheader_udiv32x_xexitx_xix_xi20_PhiReq/phi_stmt_2990/phi_stmt_2990_sources/type_cast_2993/SplitProtocol/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi20x_xpreheader_udiv32x_xexitx_xix_xi20_PhiReq/phi_stmt_2990/phi_stmt_2990_req
      -- 
    cp_element_group_1876: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1876"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1874) & cp_elements(1875);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1876), clk => clk, reset => reset); --
    end block;
    phi_stmt_2990_req_17918_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1876), ack => phi_stmt_2990_req_1); -- 
    -- CP-element group 1877 fork  transition  bypass 
    -- predecessors 1872 
    -- successors 1878 1882 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi20x_xpreheader_udiv32x_xexitx_xix_xi20_PhiReq/phi_stmt_2997/$entry
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi20x_xpreheader_udiv32x_xexitx_xix_xi20_PhiReq/phi_stmt_2997/phi_stmt_2997_sources/$entry
      -- 
    cp_elements(1877) <= cp_elements(1872);
    -- CP-element group 1878 fork  transition  bypass 
    -- predecessors 1877 
    -- successors 1879 1880 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi20x_xpreheader_udiv32x_xexitx_xix_xi20_PhiReq/phi_stmt_2997/phi_stmt_2997_sources/type_cast_3000/$entry
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi20x_xpreheader_udiv32x_xexitx_xix_xi20_PhiReq/phi_stmt_2997/phi_stmt_2997_sources/type_cast_3000/SplitProtocol/$entry
      -- 
    cp_elements(1878) <= cp_elements(1877);
    -- CP-element group 1879 transition  bypass 
    -- predecessors 1878 
    -- successors 1881 
    -- members (4) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi20x_xpreheader_udiv32x_xexitx_xix_xi20_PhiReq/phi_stmt_2997/phi_stmt_2997_sources/type_cast_3000/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi20x_xpreheader_udiv32x_xexitx_xix_xi20_PhiReq/phi_stmt_2997/phi_stmt_2997_sources/type_cast_3000/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi20x_xpreheader_udiv32x_xexitx_xix_xi20_PhiReq/phi_stmt_2997/phi_stmt_2997_sources/type_cast_3000/SplitProtocol/Sample/rr
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi20x_xpreheader_udiv32x_xexitx_xix_xi20_PhiReq/phi_stmt_2997/phi_stmt_2997_sources/type_cast_3000/SplitProtocol/Sample/ra
      -- 
    cp_elements(1879) <= cp_elements(1878);
    -- CP-element group 1880 transition  bypass 
    -- predecessors 1878 
    -- successors 1881 
    -- members (4) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi20x_xpreheader_udiv32x_xexitx_xix_xi20_PhiReq/phi_stmt_2997/phi_stmt_2997_sources/type_cast_3000/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi20x_xpreheader_udiv32x_xexitx_xix_xi20_PhiReq/phi_stmt_2997/phi_stmt_2997_sources/type_cast_3000/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi20x_xpreheader_udiv32x_xexitx_xix_xi20_PhiReq/phi_stmt_2997/phi_stmt_2997_sources/type_cast_3000/SplitProtocol/Update/cr
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi20x_xpreheader_udiv32x_xexitx_xix_xi20_PhiReq/phi_stmt_2997/phi_stmt_2997_sources/type_cast_3000/SplitProtocol/Update/ca
      -- 
    cp_elements(1880) <= cp_elements(1878);
    -- CP-element group 1881 join  transition  bypass 
    -- predecessors 1879 1880 
    -- successors 1888 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi20x_xpreheader_udiv32x_xexitx_xix_xi20_PhiReq/phi_stmt_2997/phi_stmt_2997_sources/type_cast_3000/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi20x_xpreheader_udiv32x_xexitx_xix_xi20_PhiReq/phi_stmt_2997/phi_stmt_2997_sources/type_cast_3000/SplitProtocol/$exit
      -- 
    cp_element_group_1881: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1881"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1879) & cp_elements(1880);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1881), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1882 fork  transition  bypass 
    -- predecessors 1877 
    -- successors 1883 1885 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi20x_xpreheader_udiv32x_xexitx_xix_xi20_PhiReq/phi_stmt_2997/phi_stmt_2997_sources/type_cast_3002/$entry
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi20x_xpreheader_udiv32x_xexitx_xix_xi20_PhiReq/phi_stmt_2997/phi_stmt_2997_sources/type_cast_3002/SplitProtocol/$entry
      -- 
    cp_elements(1882) <= cp_elements(1877);
    -- CP-element group 1883 transition  output  bypass 
    -- predecessors 1882 
    -- successors 1884 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi20x_xpreheader_udiv32x_xexitx_xix_xi20_PhiReq/phi_stmt_2997/phi_stmt_2997_sources/type_cast_3002/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi20x_xpreheader_udiv32x_xexitx_xix_xi20_PhiReq/phi_stmt_2997/phi_stmt_2997_sources/type_cast_3002/SplitProtocol/Sample/rr
      -- 
    cp_elements(1883) <= cp_elements(1882);
    rr_17950_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1883), ack => type_cast_3002_inst_req_0); -- 
    -- CP-element group 1884 transition  input  bypass 
    -- predecessors 1883 
    -- successors 1887 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi20x_xpreheader_udiv32x_xexitx_xix_xi20_PhiReq/phi_stmt_2997/phi_stmt_2997_sources/type_cast_3002/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi20x_xpreheader_udiv32x_xexitx_xix_xi20_PhiReq/phi_stmt_2997/phi_stmt_2997_sources/type_cast_3002/SplitProtocol/Sample/ra
      -- 
    ra_17951_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3002_inst_ack_0, ack => cp_elements(1884)); -- 
    -- CP-element group 1885 transition  output  bypass 
    -- predecessors 1882 
    -- successors 1886 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi20x_xpreheader_udiv32x_xexitx_xix_xi20_PhiReq/phi_stmt_2997/phi_stmt_2997_sources/type_cast_3002/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi20x_xpreheader_udiv32x_xexitx_xix_xi20_PhiReq/phi_stmt_2997/phi_stmt_2997_sources/type_cast_3002/SplitProtocol/Update/cr
      -- 
    cp_elements(1885) <= cp_elements(1882);
    cr_17955_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1885), ack => type_cast_3002_inst_req_1); -- 
    -- CP-element group 1886 transition  input  bypass 
    -- predecessors 1885 
    -- successors 1887 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi20x_xpreheader_udiv32x_xexitx_xix_xi20_PhiReq/phi_stmt_2997/phi_stmt_2997_sources/type_cast_3002/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi20x_xpreheader_udiv32x_xexitx_xix_xi20_PhiReq/phi_stmt_2997/phi_stmt_2997_sources/type_cast_3002/SplitProtocol/Update/ca
      -- 
    ca_17956_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3002_inst_ack_1, ack => cp_elements(1886)); -- 
    -- CP-element group 1887 join  transition  bypass 
    -- predecessors 1884 1886 
    -- successors 1888 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi20x_xpreheader_udiv32x_xexitx_xix_xi20_PhiReq/phi_stmt_2997/phi_stmt_2997_sources/type_cast_3002/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi20x_xpreheader_udiv32x_xexitx_xix_xi20_PhiReq/phi_stmt_2997/phi_stmt_2997_sources/type_cast_3002/SplitProtocol/$exit
      -- 
    cp_element_group_1887: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1887"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1884) & cp_elements(1886);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1887), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1888 join  transition  output  bypass 
    -- predecessors 1881 1887 
    -- successors 1889 
    -- members (3) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi20x_xpreheader_udiv32x_xexitx_xix_xi20_PhiReq/phi_stmt_2997/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi20x_xpreheader_udiv32x_xexitx_xix_xi20_PhiReq/phi_stmt_2997/phi_stmt_2997_sources/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi20x_xpreheader_udiv32x_xexitx_xix_xi20_PhiReq/phi_stmt_2997/phi_stmt_2997_req
      -- 
    cp_element_group_1888: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1888"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1881) & cp_elements(1887);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1888), clk => clk, reset => reset); --
    end block;
    phi_stmt_2997_req_17957_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1888), ack => phi_stmt_2997_req_1); -- 
    -- CP-element group 1889 join  transition  bypass 
    -- predecessors 1876 1888 
    -- successors 1890 
    -- members (1) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi20x_xpreheader_udiv32x_xexitx_xix_xi20_PhiReq/$exit
      -- 
    cp_element_group_1889: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1889"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1876) & cp_elements(1888);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1889), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1890 merge  place  bypass 
    -- predecessors 1871 1889 
    -- successors 1891 
    -- members (1) 
      -- 	branch_block_stmt_2042/merge_stmt_2989_PhiReqMerge
      -- 
    cp_elements(1890) <= OrReduce(cp_elements(1871) & cp_elements(1889));
    -- CP-element group 1891 fork  transition  bypass 
    -- predecessors 1890 
    -- successors 1892 1893 
    -- members (1) 
      -- 	branch_block_stmt_2042/merge_stmt_2989_PhiAck/$entry
      -- 
    cp_elements(1891) <= cp_elements(1890);
    -- CP-element group 1892 transition  input  bypass 
    -- predecessors 1891 
    -- successors 1894 
    -- members (1) 
      -- 	branch_block_stmt_2042/merge_stmt_2989_PhiAck/phi_stmt_2990_ack
      -- 
    phi_stmt_2990_ack_17962_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2990_ack_0, ack => cp_elements(1892)); -- 
    -- CP-element group 1893 transition  input  bypass 
    -- predecessors 1891 
    -- successors 1894 
    -- members (1) 
      -- 	branch_block_stmt_2042/merge_stmt_2989_PhiAck/phi_stmt_2997_ack
      -- 
    phi_stmt_2997_ack_17963_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2997_ack_0, ack => cp_elements(1893)); -- 
    -- CP-element group 1894 join  transition  bypass 
    -- predecessors 1892 1893 
    -- successors 39 
    -- members (1) 
      -- 	branch_block_stmt_2042/merge_stmt_2989_PhiAck/$exit
      -- 
    cp_element_group_1894: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1894"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1892) & cp_elements(1893);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1894), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1895 fork  transition  bypass 
    -- predecessors 683 
    -- successors 1896 1902 
    -- members (1) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi20_udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi24_PhiReq/$entry
      -- 
    cp_elements(1895) <= cp_elements(683);
    -- CP-element group 1896 fork  transition  bypass 
    -- predecessors 1895 
    -- successors 1897 1899 
    -- members (4) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi20_udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi24_PhiReq/phi_stmt_3048/$entry
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi20_udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi24_PhiReq/phi_stmt_3048/phi_stmt_3048_sources/$entry
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi20_udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi24_PhiReq/phi_stmt_3048/phi_stmt_3048_sources/type_cast_3051/$entry
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi20_udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi24_PhiReq/phi_stmt_3048/phi_stmt_3048_sources/type_cast_3051/SplitProtocol/$entry
      -- 
    cp_elements(1896) <= cp_elements(1895);
    -- CP-element group 1897 transition  output  bypass 
    -- predecessors 1896 
    -- successors 1898 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi20_udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi24_PhiReq/phi_stmt_3048/phi_stmt_3048_sources/type_cast_3051/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi20_udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi24_PhiReq/phi_stmt_3048/phi_stmt_3048_sources/type_cast_3051/SplitProtocol/Sample/rr
      -- 
    cp_elements(1897) <= cp_elements(1896);
    rr_17986_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1897), ack => type_cast_3051_inst_req_0); -- 
    -- CP-element group 1898 transition  input  bypass 
    -- predecessors 1897 
    -- successors 1901 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi20_udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi24_PhiReq/phi_stmt_3048/phi_stmt_3048_sources/type_cast_3051/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi20_udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi24_PhiReq/phi_stmt_3048/phi_stmt_3048_sources/type_cast_3051/SplitProtocol/Sample/ra
      -- 
    ra_17987_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3051_inst_ack_0, ack => cp_elements(1898)); -- 
    -- CP-element group 1899 transition  output  bypass 
    -- predecessors 1896 
    -- successors 1900 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi20_udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi24_PhiReq/phi_stmt_3048/phi_stmt_3048_sources/type_cast_3051/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi20_udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi24_PhiReq/phi_stmt_3048/phi_stmt_3048_sources/type_cast_3051/SplitProtocol/Update/cr
      -- 
    cp_elements(1899) <= cp_elements(1896);
    cr_17991_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1899), ack => type_cast_3051_inst_req_1); -- 
    -- CP-element group 1900 transition  input  bypass 
    -- predecessors 1899 
    -- successors 1901 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi20_udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi24_PhiReq/phi_stmt_3048/phi_stmt_3048_sources/type_cast_3051/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi20_udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi24_PhiReq/phi_stmt_3048/phi_stmt_3048_sources/type_cast_3051/SplitProtocol/Update/ca
      -- 
    ca_17992_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3051_inst_ack_1, ack => cp_elements(1900)); -- 
    -- CP-element group 1901 join  transition  output  bypass 
    -- predecessors 1898 1900 
    -- successors 1908 
    -- members (5) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi20_udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi24_PhiReq/phi_stmt_3048/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi20_udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi24_PhiReq/phi_stmt_3048/phi_stmt_3048_sources/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi20_udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi24_PhiReq/phi_stmt_3048/phi_stmt_3048_sources/type_cast_3051/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi20_udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi24_PhiReq/phi_stmt_3048/phi_stmt_3048_sources/type_cast_3051/SplitProtocol/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi20_udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi24_PhiReq/phi_stmt_3048/phi_stmt_3048_req
      -- 
    cp_element_group_1901: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1901"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1898) & cp_elements(1900);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1901), clk => clk, reset => reset); --
    end block;
    phi_stmt_3048_req_17993_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1901), ack => phi_stmt_3048_req_0); -- 
    -- CP-element group 1902 fork  transition  bypass 
    -- predecessors 1895 
    -- successors 1903 1905 
    -- members (4) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi20_udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi24_PhiReq/phi_stmt_3052/$entry
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi20_udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi24_PhiReq/phi_stmt_3052/phi_stmt_3052_sources/$entry
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi20_udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi24_PhiReq/phi_stmt_3052/phi_stmt_3052_sources/type_cast_3055/$entry
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi20_udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi24_PhiReq/phi_stmt_3052/phi_stmt_3052_sources/type_cast_3055/SplitProtocol/$entry
      -- 
    cp_elements(1902) <= cp_elements(1895);
    -- CP-element group 1903 transition  output  bypass 
    -- predecessors 1902 
    -- successors 1904 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi20_udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi24_PhiReq/phi_stmt_3052/phi_stmt_3052_sources/type_cast_3055/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi20_udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi24_PhiReq/phi_stmt_3052/phi_stmt_3052_sources/type_cast_3055/SplitProtocol/Sample/rr
      -- 
    cp_elements(1903) <= cp_elements(1902);
    rr_18009_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1903), ack => type_cast_3055_inst_req_0); -- 
    -- CP-element group 1904 transition  input  bypass 
    -- predecessors 1903 
    -- successors 1907 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi20_udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi24_PhiReq/phi_stmt_3052/phi_stmt_3052_sources/type_cast_3055/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi20_udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi24_PhiReq/phi_stmt_3052/phi_stmt_3052_sources/type_cast_3055/SplitProtocol/Sample/ra
      -- 
    ra_18010_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3055_inst_ack_0, ack => cp_elements(1904)); -- 
    -- CP-element group 1905 transition  output  bypass 
    -- predecessors 1902 
    -- successors 1906 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi20_udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi24_PhiReq/phi_stmt_3052/phi_stmt_3052_sources/type_cast_3055/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi20_udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi24_PhiReq/phi_stmt_3052/phi_stmt_3052_sources/type_cast_3055/SplitProtocol/Update/cr
      -- 
    cp_elements(1905) <= cp_elements(1902);
    cr_18014_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1905), ack => type_cast_3055_inst_req_1); -- 
    -- CP-element group 1906 transition  input  bypass 
    -- predecessors 1905 
    -- successors 1907 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi20_udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi24_PhiReq/phi_stmt_3052/phi_stmt_3052_sources/type_cast_3055/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi20_udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi24_PhiReq/phi_stmt_3052/phi_stmt_3052_sources/type_cast_3055/SplitProtocol/Update/ca
      -- 
    ca_18015_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3055_inst_ack_1, ack => cp_elements(1906)); -- 
    -- CP-element group 1907 join  transition  output  bypass 
    -- predecessors 1904 1906 
    -- successors 1908 
    -- members (5) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi20_udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi24_PhiReq/phi_stmt_3052/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi20_udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi24_PhiReq/phi_stmt_3052/phi_stmt_3052_sources/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi20_udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi24_PhiReq/phi_stmt_3052/phi_stmt_3052_sources/type_cast_3055/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi20_udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi24_PhiReq/phi_stmt_3052/phi_stmt_3052_sources/type_cast_3055/SplitProtocol/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi20_udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi24_PhiReq/phi_stmt_3052/phi_stmt_3052_req
      -- 
    cp_element_group_1907: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1907"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1904) & cp_elements(1906);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1907), clk => clk, reset => reset); --
    end block;
    phi_stmt_3052_req_18016_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1907), ack => phi_stmt_3052_req_0); -- 
    -- CP-element group 1908 join  transition  bypass 
    -- predecessors 1901 1907 
    -- successors 1909 
    -- members (1) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi20_udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi24_PhiReq/$exit
      -- 
    cp_element_group_1908: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1908"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1901) & cp_elements(1907);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1908), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1909 place  bypass 
    -- predecessors 1908 
    -- successors 1910 
    -- members (1) 
      -- 	branch_block_stmt_2042/merge_stmt_3047_PhiReqMerge
      -- 
    cp_elements(1909) <= cp_elements(1908);
    -- CP-element group 1910 fork  transition  bypass 
    -- predecessors 1909 
    -- successors 1911 1912 
    -- members (1) 
      -- 	branch_block_stmt_2042/merge_stmt_3047_PhiAck/$entry
      -- 
    cp_elements(1910) <= cp_elements(1909);
    -- CP-element group 1911 transition  input  bypass 
    -- predecessors 1910 
    -- successors 1913 
    -- members (1) 
      -- 	branch_block_stmt_2042/merge_stmt_3047_PhiAck/phi_stmt_3048_ack
      -- 
    phi_stmt_3048_ack_18021_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_3048_ack_0, ack => cp_elements(1911)); -- 
    -- CP-element group 1912 transition  input  bypass 
    -- predecessors 1910 
    -- successors 1913 
    -- members (1) 
      -- 	branch_block_stmt_2042/merge_stmt_3047_PhiAck/phi_stmt_3052_ack
      -- 
    phi_stmt_3052_ack_18022_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_3052_ack_0, ack => cp_elements(1912)); -- 
    -- CP-element group 1913 join  transition  bypass 
    -- predecessors 1911 1912 
    -- successors 41 
    -- members (1) 
      -- 	branch_block_stmt_2042/merge_stmt_3047_PhiAck/$exit
      -- 
    cp_element_group_1913: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1913"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1911) & cp_elements(1912);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1913), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1914 fork  transition  bypass 
    -- predecessors 649 
    -- successors 1915 1927 
    -- members (1) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xpreheaderx_xix_xi16_xx_xcritedgex_xix_xi28_PhiReq/$entry
      -- 
    cp_elements(1914) <= cp_elements(649);
    -- CP-element group 1915 fork  transition  bypass 
    -- predecessors 1914 
    -- successors 1916 1920 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xpreheaderx_xix_xi16_xx_xcritedgex_xix_xi28_PhiReq/phi_stmt_3075/$entry
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xpreheaderx_xix_xi16_xx_xcritedgex_xix_xi28_PhiReq/phi_stmt_3075/phi_stmt_3075_sources/$entry
      -- 
    cp_elements(1915) <= cp_elements(1914);
    -- CP-element group 1916 fork  transition  bypass 
    -- predecessors 1915 
    -- successors 1917 1918 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xpreheaderx_xix_xi16_xx_xcritedgex_xix_xi28_PhiReq/phi_stmt_3075/phi_stmt_3075_sources/type_cast_3078/$entry
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xpreheaderx_xix_xi16_xx_xcritedgex_xix_xi28_PhiReq/phi_stmt_3075/phi_stmt_3075_sources/type_cast_3078/SplitProtocol/$entry
      -- 
    cp_elements(1916) <= cp_elements(1915);
    -- CP-element group 1917 transition  bypass 
    -- predecessors 1916 
    -- successors 1919 
    -- members (4) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xpreheaderx_xix_xi16_xx_xcritedgex_xix_xi28_PhiReq/phi_stmt_3075/phi_stmt_3075_sources/type_cast_3078/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xpreheaderx_xix_xi16_xx_xcritedgex_xix_xi28_PhiReq/phi_stmt_3075/phi_stmt_3075_sources/type_cast_3078/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xpreheaderx_xix_xi16_xx_xcritedgex_xix_xi28_PhiReq/phi_stmt_3075/phi_stmt_3075_sources/type_cast_3078/SplitProtocol/Sample/rr
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xpreheaderx_xix_xi16_xx_xcritedgex_xix_xi28_PhiReq/phi_stmt_3075/phi_stmt_3075_sources/type_cast_3078/SplitProtocol/Sample/ra
      -- 
    cp_elements(1917) <= cp_elements(1916);
    -- CP-element group 1918 transition  bypass 
    -- predecessors 1916 
    -- successors 1919 
    -- members (4) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xpreheaderx_xix_xi16_xx_xcritedgex_xix_xi28_PhiReq/phi_stmt_3075/phi_stmt_3075_sources/type_cast_3078/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xpreheaderx_xix_xi16_xx_xcritedgex_xix_xi28_PhiReq/phi_stmt_3075/phi_stmt_3075_sources/type_cast_3078/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xpreheaderx_xix_xi16_xx_xcritedgex_xix_xi28_PhiReq/phi_stmt_3075/phi_stmt_3075_sources/type_cast_3078/SplitProtocol/Update/cr
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xpreheaderx_xix_xi16_xx_xcritedgex_xix_xi28_PhiReq/phi_stmt_3075/phi_stmt_3075_sources/type_cast_3078/SplitProtocol/Update/ca
      -- 
    cp_elements(1918) <= cp_elements(1916);
    -- CP-element group 1919 join  transition  bypass 
    -- predecessors 1917 1918 
    -- successors 1926 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xpreheaderx_xix_xi16_xx_xcritedgex_xix_xi28_PhiReq/phi_stmt_3075/phi_stmt_3075_sources/type_cast_3078/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xpreheaderx_xix_xi16_xx_xcritedgex_xix_xi28_PhiReq/phi_stmt_3075/phi_stmt_3075_sources/type_cast_3078/SplitProtocol/$exit
      -- 
    cp_element_group_1919: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1919"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1917) & cp_elements(1918);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1919), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1920 fork  transition  bypass 
    -- predecessors 1915 
    -- successors 1921 1923 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xpreheaderx_xix_xi16_xx_xcritedgex_xix_xi28_PhiReq/phi_stmt_3075/phi_stmt_3075_sources/type_cast_3080/$entry
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xpreheaderx_xix_xi16_xx_xcritedgex_xix_xi28_PhiReq/phi_stmt_3075/phi_stmt_3075_sources/type_cast_3080/SplitProtocol/$entry
      -- 
    cp_elements(1920) <= cp_elements(1915);
    -- CP-element group 1921 transition  output  bypass 
    -- predecessors 1920 
    -- successors 1922 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xpreheaderx_xix_xi16_xx_xcritedgex_xix_xi28_PhiReq/phi_stmt_3075/phi_stmt_3075_sources/type_cast_3080/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xpreheaderx_xix_xi16_xx_xcritedgex_xix_xi28_PhiReq/phi_stmt_3075/phi_stmt_3075_sources/type_cast_3080/SplitProtocol/Sample/rr
      -- 
    cp_elements(1921) <= cp_elements(1920);
    rr_18057_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1921), ack => type_cast_3080_inst_req_0); -- 
    -- CP-element group 1922 transition  input  bypass 
    -- predecessors 1921 
    -- successors 1925 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xpreheaderx_xix_xi16_xx_xcritedgex_xix_xi28_PhiReq/phi_stmt_3075/phi_stmt_3075_sources/type_cast_3080/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xpreheaderx_xix_xi16_xx_xcritedgex_xix_xi28_PhiReq/phi_stmt_3075/phi_stmt_3075_sources/type_cast_3080/SplitProtocol/Sample/ra
      -- 
    ra_18058_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3080_inst_ack_0, ack => cp_elements(1922)); -- 
    -- CP-element group 1923 transition  output  bypass 
    -- predecessors 1920 
    -- successors 1924 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xpreheaderx_xix_xi16_xx_xcritedgex_xix_xi28_PhiReq/phi_stmt_3075/phi_stmt_3075_sources/type_cast_3080/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xpreheaderx_xix_xi16_xx_xcritedgex_xix_xi28_PhiReq/phi_stmt_3075/phi_stmt_3075_sources/type_cast_3080/SplitProtocol/Update/cr
      -- 
    cp_elements(1923) <= cp_elements(1920);
    cr_18062_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1923), ack => type_cast_3080_inst_req_1); -- 
    -- CP-element group 1924 transition  input  bypass 
    -- predecessors 1923 
    -- successors 1925 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xpreheaderx_xix_xi16_xx_xcritedgex_xix_xi28_PhiReq/phi_stmt_3075/phi_stmt_3075_sources/type_cast_3080/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xpreheaderx_xix_xi16_xx_xcritedgex_xix_xi28_PhiReq/phi_stmt_3075/phi_stmt_3075_sources/type_cast_3080/SplitProtocol/Update/ca
      -- 
    ca_18063_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3080_inst_ack_1, ack => cp_elements(1924)); -- 
    -- CP-element group 1925 join  transition  bypass 
    -- predecessors 1922 1924 
    -- successors 1926 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xpreheaderx_xix_xi16_xx_xcritedgex_xix_xi28_PhiReq/phi_stmt_3075/phi_stmt_3075_sources/type_cast_3080/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xpreheaderx_xix_xi16_xx_xcritedgex_xix_xi28_PhiReq/phi_stmt_3075/phi_stmt_3075_sources/type_cast_3080/SplitProtocol/$exit
      -- 
    cp_element_group_1925: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1925"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1922) & cp_elements(1924);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1925), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1926 join  transition  output  bypass 
    -- predecessors 1919 1925 
    -- successors 1939 
    -- members (3) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xpreheaderx_xix_xi16_xx_xcritedgex_xix_xi28_PhiReq/phi_stmt_3075/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xpreheaderx_xix_xi16_xx_xcritedgex_xix_xi28_PhiReq/phi_stmt_3075/phi_stmt_3075_sources/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xpreheaderx_xix_xi16_xx_xcritedgex_xix_xi28_PhiReq/phi_stmt_3075/phi_stmt_3075_req
      -- 
    cp_element_group_1926: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1926"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1919) & cp_elements(1925);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1926), clk => clk, reset => reset); --
    end block;
    phi_stmt_3075_req_18064_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1926), ack => phi_stmt_3075_req_1); -- 
    -- CP-element group 1927 fork  transition  bypass 
    -- predecessors 1914 
    -- successors 1928 1932 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xpreheaderx_xix_xi16_xx_xcritedgex_xix_xi28_PhiReq/phi_stmt_3081/$entry
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xpreheaderx_xix_xi16_xx_xcritedgex_xix_xi28_PhiReq/phi_stmt_3081/phi_stmt_3081_sources/$entry
      -- 
    cp_elements(1927) <= cp_elements(1914);
    -- CP-element group 1928 fork  transition  bypass 
    -- predecessors 1927 
    -- successors 1929 1930 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xpreheaderx_xix_xi16_xx_xcritedgex_xix_xi28_PhiReq/phi_stmt_3081/phi_stmt_3081_sources/type_cast_3084/$entry
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xpreheaderx_xix_xi16_xx_xcritedgex_xix_xi28_PhiReq/phi_stmt_3081/phi_stmt_3081_sources/type_cast_3084/SplitProtocol/$entry
      -- 
    cp_elements(1928) <= cp_elements(1927);
    -- CP-element group 1929 transition  bypass 
    -- predecessors 1928 
    -- successors 1931 
    -- members (4) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xpreheaderx_xix_xi16_xx_xcritedgex_xix_xi28_PhiReq/phi_stmt_3081/phi_stmt_3081_sources/type_cast_3084/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xpreheaderx_xix_xi16_xx_xcritedgex_xix_xi28_PhiReq/phi_stmt_3081/phi_stmt_3081_sources/type_cast_3084/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xpreheaderx_xix_xi16_xx_xcritedgex_xix_xi28_PhiReq/phi_stmt_3081/phi_stmt_3081_sources/type_cast_3084/SplitProtocol/Sample/rr
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xpreheaderx_xix_xi16_xx_xcritedgex_xix_xi28_PhiReq/phi_stmt_3081/phi_stmt_3081_sources/type_cast_3084/SplitProtocol/Sample/ra
      -- 
    cp_elements(1929) <= cp_elements(1928);
    -- CP-element group 1930 transition  bypass 
    -- predecessors 1928 
    -- successors 1931 
    -- members (4) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xpreheaderx_xix_xi16_xx_xcritedgex_xix_xi28_PhiReq/phi_stmt_3081/phi_stmt_3081_sources/type_cast_3084/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xpreheaderx_xix_xi16_xx_xcritedgex_xix_xi28_PhiReq/phi_stmt_3081/phi_stmt_3081_sources/type_cast_3084/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xpreheaderx_xix_xi16_xx_xcritedgex_xix_xi28_PhiReq/phi_stmt_3081/phi_stmt_3081_sources/type_cast_3084/SplitProtocol/Update/cr
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xpreheaderx_xix_xi16_xx_xcritedgex_xix_xi28_PhiReq/phi_stmt_3081/phi_stmt_3081_sources/type_cast_3084/SplitProtocol/Update/ca
      -- 
    cp_elements(1930) <= cp_elements(1928);
    -- CP-element group 1931 join  transition  bypass 
    -- predecessors 1929 1930 
    -- successors 1938 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xpreheaderx_xix_xi16_xx_xcritedgex_xix_xi28_PhiReq/phi_stmt_3081/phi_stmt_3081_sources/type_cast_3084/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xpreheaderx_xix_xi16_xx_xcritedgex_xix_xi28_PhiReq/phi_stmt_3081/phi_stmt_3081_sources/type_cast_3084/SplitProtocol/$exit
      -- 
    cp_element_group_1931: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1931"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1929) & cp_elements(1930);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1931), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1932 fork  transition  bypass 
    -- predecessors 1927 
    -- successors 1933 1935 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xpreheaderx_xix_xi16_xx_xcritedgex_xix_xi28_PhiReq/phi_stmt_3081/phi_stmt_3081_sources/type_cast_3086/$entry
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xpreheaderx_xix_xi16_xx_xcritedgex_xix_xi28_PhiReq/phi_stmt_3081/phi_stmt_3081_sources/type_cast_3086/SplitProtocol/$entry
      -- 
    cp_elements(1932) <= cp_elements(1927);
    -- CP-element group 1933 transition  output  bypass 
    -- predecessors 1932 
    -- successors 1934 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xpreheaderx_xix_xi16_xx_xcritedgex_xix_xi28_PhiReq/phi_stmt_3081/phi_stmt_3081_sources/type_cast_3086/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xpreheaderx_xix_xi16_xx_xcritedgex_xix_xi28_PhiReq/phi_stmt_3081/phi_stmt_3081_sources/type_cast_3086/SplitProtocol/Sample/rr
      -- 
    cp_elements(1933) <= cp_elements(1932);
    rr_18096_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1933), ack => type_cast_3086_inst_req_0); -- 
    -- CP-element group 1934 transition  input  bypass 
    -- predecessors 1933 
    -- successors 1937 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xpreheaderx_xix_xi16_xx_xcritedgex_xix_xi28_PhiReq/phi_stmt_3081/phi_stmt_3081_sources/type_cast_3086/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xpreheaderx_xix_xi16_xx_xcritedgex_xix_xi28_PhiReq/phi_stmt_3081/phi_stmt_3081_sources/type_cast_3086/SplitProtocol/Sample/ra
      -- 
    ra_18097_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3086_inst_ack_0, ack => cp_elements(1934)); -- 
    -- CP-element group 1935 transition  output  bypass 
    -- predecessors 1932 
    -- successors 1936 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xpreheaderx_xix_xi16_xx_xcritedgex_xix_xi28_PhiReq/phi_stmt_3081/phi_stmt_3081_sources/type_cast_3086/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xpreheaderx_xix_xi16_xx_xcritedgex_xix_xi28_PhiReq/phi_stmt_3081/phi_stmt_3081_sources/type_cast_3086/SplitProtocol/Update/cr
      -- 
    cp_elements(1935) <= cp_elements(1932);
    cr_18101_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1935), ack => type_cast_3086_inst_req_1); -- 
    -- CP-element group 1936 transition  input  bypass 
    -- predecessors 1935 
    -- successors 1937 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xpreheaderx_xix_xi16_xx_xcritedgex_xix_xi28_PhiReq/phi_stmt_3081/phi_stmt_3081_sources/type_cast_3086/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xpreheaderx_xix_xi16_xx_xcritedgex_xix_xi28_PhiReq/phi_stmt_3081/phi_stmt_3081_sources/type_cast_3086/SplitProtocol/Update/ca
      -- 
    ca_18102_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3086_inst_ack_1, ack => cp_elements(1936)); -- 
    -- CP-element group 1937 join  transition  bypass 
    -- predecessors 1934 1936 
    -- successors 1938 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xpreheaderx_xix_xi16_xx_xcritedgex_xix_xi28_PhiReq/phi_stmt_3081/phi_stmt_3081_sources/type_cast_3086/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xpreheaderx_xix_xi16_xx_xcritedgex_xix_xi28_PhiReq/phi_stmt_3081/phi_stmt_3081_sources/type_cast_3086/SplitProtocol/$exit
      -- 
    cp_element_group_1937: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1937"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1934) & cp_elements(1936);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1937), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1938 join  transition  output  bypass 
    -- predecessors 1931 1937 
    -- successors 1939 
    -- members (3) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xpreheaderx_xix_xi16_xx_xcritedgex_xix_xi28_PhiReq/phi_stmt_3081/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xpreheaderx_xix_xi16_xx_xcritedgex_xix_xi28_PhiReq/phi_stmt_3081/phi_stmt_3081_sources/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xpreheaderx_xix_xi16_xx_xcritedgex_xix_xi28_PhiReq/phi_stmt_3081/phi_stmt_3081_req
      -- 
    cp_element_group_1938: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1938"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1931) & cp_elements(1937);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1938), clk => clk, reset => reset); --
    end block;
    phi_stmt_3081_req_18103_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1938), ack => phi_stmt_3081_req_1); -- 
    -- CP-element group 1939 join  transition  bypass 
    -- predecessors 1926 1938 
    -- successors 1966 
    -- members (1) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xpreheaderx_xix_xi16_xx_xcritedgex_xix_xi28_PhiReq/$exit
      -- 
    cp_element_group_1939: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1939"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1926) & cp_elements(1938);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1939), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1940 fork  transition  bypass 
    -- predecessors 698 
    -- successors 1941 1953 
    -- members (1) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi24_xx_xcritedgex_xix_xi28_PhiReq/$entry
      -- 
    cp_elements(1940) <= cp_elements(698);
    -- CP-element group 1941 fork  transition  bypass 
    -- predecessors 1940 
    -- successors 1942 1948 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi24_xx_xcritedgex_xix_xi28_PhiReq/phi_stmt_3075/$entry
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi24_xx_xcritedgex_xix_xi28_PhiReq/phi_stmt_3075/phi_stmt_3075_sources/$entry
      -- 
    cp_elements(1941) <= cp_elements(1940);
    -- CP-element group 1942 fork  transition  bypass 
    -- predecessors 1941 
    -- successors 1943 1945 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi24_xx_xcritedgex_xix_xi28_PhiReq/phi_stmt_3075/phi_stmt_3075_sources/type_cast_3078/$entry
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi24_xx_xcritedgex_xix_xi28_PhiReq/phi_stmt_3075/phi_stmt_3075_sources/type_cast_3078/SplitProtocol/$entry
      -- 
    cp_elements(1942) <= cp_elements(1941);
    -- CP-element group 1943 transition  output  bypass 
    -- predecessors 1942 
    -- successors 1944 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi24_xx_xcritedgex_xix_xi28_PhiReq/phi_stmt_3075/phi_stmt_3075_sources/type_cast_3078/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi24_xx_xcritedgex_xix_xi28_PhiReq/phi_stmt_3075/phi_stmt_3075_sources/type_cast_3078/SplitProtocol/Sample/rr
      -- 
    cp_elements(1943) <= cp_elements(1942);
    rr_18122_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1943), ack => type_cast_3078_inst_req_0); -- 
    -- CP-element group 1944 transition  input  bypass 
    -- predecessors 1943 
    -- successors 1947 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi24_xx_xcritedgex_xix_xi28_PhiReq/phi_stmt_3075/phi_stmt_3075_sources/type_cast_3078/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi24_xx_xcritedgex_xix_xi28_PhiReq/phi_stmt_3075/phi_stmt_3075_sources/type_cast_3078/SplitProtocol/Sample/ra
      -- 
    ra_18123_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3078_inst_ack_0, ack => cp_elements(1944)); -- 
    -- CP-element group 1945 transition  output  bypass 
    -- predecessors 1942 
    -- successors 1946 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi24_xx_xcritedgex_xix_xi28_PhiReq/phi_stmt_3075/phi_stmt_3075_sources/type_cast_3078/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi24_xx_xcritedgex_xix_xi28_PhiReq/phi_stmt_3075/phi_stmt_3075_sources/type_cast_3078/SplitProtocol/Update/cr
      -- 
    cp_elements(1945) <= cp_elements(1942);
    cr_18127_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1945), ack => type_cast_3078_inst_req_1); -- 
    -- CP-element group 1946 transition  input  bypass 
    -- predecessors 1945 
    -- successors 1947 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi24_xx_xcritedgex_xix_xi28_PhiReq/phi_stmt_3075/phi_stmt_3075_sources/type_cast_3078/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi24_xx_xcritedgex_xix_xi28_PhiReq/phi_stmt_3075/phi_stmt_3075_sources/type_cast_3078/SplitProtocol/Update/ca
      -- 
    ca_18128_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3078_inst_ack_1, ack => cp_elements(1946)); -- 
    -- CP-element group 1947 join  transition  bypass 
    -- predecessors 1944 1946 
    -- successors 1952 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi24_xx_xcritedgex_xix_xi28_PhiReq/phi_stmt_3075/phi_stmt_3075_sources/type_cast_3078/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi24_xx_xcritedgex_xix_xi28_PhiReq/phi_stmt_3075/phi_stmt_3075_sources/type_cast_3078/SplitProtocol/$exit
      -- 
    cp_element_group_1947: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1947"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1944) & cp_elements(1946);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1947), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1948 fork  transition  bypass 
    -- predecessors 1941 
    -- successors 1949 1950 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi24_xx_xcritedgex_xix_xi28_PhiReq/phi_stmt_3075/phi_stmt_3075_sources/type_cast_3080/$entry
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi24_xx_xcritedgex_xix_xi28_PhiReq/phi_stmt_3075/phi_stmt_3075_sources/type_cast_3080/SplitProtocol/$entry
      -- 
    cp_elements(1948) <= cp_elements(1941);
    -- CP-element group 1949 transition  bypass 
    -- predecessors 1948 
    -- successors 1951 
    -- members (4) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi24_xx_xcritedgex_xix_xi28_PhiReq/phi_stmt_3075/phi_stmt_3075_sources/type_cast_3080/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi24_xx_xcritedgex_xix_xi28_PhiReq/phi_stmt_3075/phi_stmt_3075_sources/type_cast_3080/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi24_xx_xcritedgex_xix_xi28_PhiReq/phi_stmt_3075/phi_stmt_3075_sources/type_cast_3080/SplitProtocol/Sample/rr
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi24_xx_xcritedgex_xix_xi28_PhiReq/phi_stmt_3075/phi_stmt_3075_sources/type_cast_3080/SplitProtocol/Sample/ra
      -- 
    cp_elements(1949) <= cp_elements(1948);
    -- CP-element group 1950 transition  bypass 
    -- predecessors 1948 
    -- successors 1951 
    -- members (4) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi24_xx_xcritedgex_xix_xi28_PhiReq/phi_stmt_3075/phi_stmt_3075_sources/type_cast_3080/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi24_xx_xcritedgex_xix_xi28_PhiReq/phi_stmt_3075/phi_stmt_3075_sources/type_cast_3080/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi24_xx_xcritedgex_xix_xi28_PhiReq/phi_stmt_3075/phi_stmt_3075_sources/type_cast_3080/SplitProtocol/Update/cr
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi24_xx_xcritedgex_xix_xi28_PhiReq/phi_stmt_3075/phi_stmt_3075_sources/type_cast_3080/SplitProtocol/Update/ca
      -- 
    cp_elements(1950) <= cp_elements(1948);
    -- CP-element group 1951 join  transition  bypass 
    -- predecessors 1949 1950 
    -- successors 1952 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi24_xx_xcritedgex_xix_xi28_PhiReq/phi_stmt_3075/phi_stmt_3075_sources/type_cast_3080/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi24_xx_xcritedgex_xix_xi28_PhiReq/phi_stmt_3075/phi_stmt_3075_sources/type_cast_3080/SplitProtocol/$exit
      -- 
    cp_element_group_1951: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1951"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1949) & cp_elements(1950);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1951), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1952 join  transition  output  bypass 
    -- predecessors 1947 1951 
    -- successors 1965 
    -- members (3) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi24_xx_xcritedgex_xix_xi28_PhiReq/phi_stmt_3075/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi24_xx_xcritedgex_xix_xi28_PhiReq/phi_stmt_3075/phi_stmt_3075_sources/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi24_xx_xcritedgex_xix_xi28_PhiReq/phi_stmt_3075/phi_stmt_3075_req
      -- 
    cp_element_group_1952: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1952"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1947) & cp_elements(1951);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1952), clk => clk, reset => reset); --
    end block;
    phi_stmt_3075_req_18145_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1952), ack => phi_stmt_3075_req_0); -- 
    -- CP-element group 1953 fork  transition  bypass 
    -- predecessors 1940 
    -- successors 1954 1960 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi24_xx_xcritedgex_xix_xi28_PhiReq/phi_stmt_3081/$entry
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi24_xx_xcritedgex_xix_xi28_PhiReq/phi_stmt_3081/phi_stmt_3081_sources/$entry
      -- 
    cp_elements(1953) <= cp_elements(1940);
    -- CP-element group 1954 fork  transition  bypass 
    -- predecessors 1953 
    -- successors 1955 1957 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi24_xx_xcritedgex_xix_xi28_PhiReq/phi_stmt_3081/phi_stmt_3081_sources/type_cast_3084/$entry
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi24_xx_xcritedgex_xix_xi28_PhiReq/phi_stmt_3081/phi_stmt_3081_sources/type_cast_3084/SplitProtocol/$entry
      -- 
    cp_elements(1954) <= cp_elements(1953);
    -- CP-element group 1955 transition  output  bypass 
    -- predecessors 1954 
    -- successors 1956 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi24_xx_xcritedgex_xix_xi28_PhiReq/phi_stmt_3081/phi_stmt_3081_sources/type_cast_3084/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi24_xx_xcritedgex_xix_xi28_PhiReq/phi_stmt_3081/phi_stmt_3081_sources/type_cast_3084/SplitProtocol/Sample/rr
      -- 
    cp_elements(1955) <= cp_elements(1954);
    rr_18161_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1955), ack => type_cast_3084_inst_req_0); -- 
    -- CP-element group 1956 transition  input  bypass 
    -- predecessors 1955 
    -- successors 1959 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi24_xx_xcritedgex_xix_xi28_PhiReq/phi_stmt_3081/phi_stmt_3081_sources/type_cast_3084/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi24_xx_xcritedgex_xix_xi28_PhiReq/phi_stmt_3081/phi_stmt_3081_sources/type_cast_3084/SplitProtocol/Sample/ra
      -- 
    ra_18162_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3084_inst_ack_0, ack => cp_elements(1956)); -- 
    -- CP-element group 1957 transition  output  bypass 
    -- predecessors 1954 
    -- successors 1958 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi24_xx_xcritedgex_xix_xi28_PhiReq/phi_stmt_3081/phi_stmt_3081_sources/type_cast_3084/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi24_xx_xcritedgex_xix_xi28_PhiReq/phi_stmt_3081/phi_stmt_3081_sources/type_cast_3084/SplitProtocol/Update/cr
      -- 
    cp_elements(1957) <= cp_elements(1954);
    cr_18166_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1957), ack => type_cast_3084_inst_req_1); -- 
    -- CP-element group 1958 transition  input  bypass 
    -- predecessors 1957 
    -- successors 1959 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi24_xx_xcritedgex_xix_xi28_PhiReq/phi_stmt_3081/phi_stmt_3081_sources/type_cast_3084/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi24_xx_xcritedgex_xix_xi28_PhiReq/phi_stmt_3081/phi_stmt_3081_sources/type_cast_3084/SplitProtocol/Update/ca
      -- 
    ca_18167_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3084_inst_ack_1, ack => cp_elements(1958)); -- 
    -- CP-element group 1959 join  transition  bypass 
    -- predecessors 1956 1958 
    -- successors 1964 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi24_xx_xcritedgex_xix_xi28_PhiReq/phi_stmt_3081/phi_stmt_3081_sources/type_cast_3084/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi24_xx_xcritedgex_xix_xi28_PhiReq/phi_stmt_3081/phi_stmt_3081_sources/type_cast_3084/SplitProtocol/$exit
      -- 
    cp_element_group_1959: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1959"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1956) & cp_elements(1958);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1959), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1960 fork  transition  bypass 
    -- predecessors 1953 
    -- successors 1961 1962 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi24_xx_xcritedgex_xix_xi28_PhiReq/phi_stmt_3081/phi_stmt_3081_sources/type_cast_3086/$entry
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi24_xx_xcritedgex_xix_xi28_PhiReq/phi_stmt_3081/phi_stmt_3081_sources/type_cast_3086/SplitProtocol/$entry
      -- 
    cp_elements(1960) <= cp_elements(1953);
    -- CP-element group 1961 transition  bypass 
    -- predecessors 1960 
    -- successors 1963 
    -- members (4) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi24_xx_xcritedgex_xix_xi28_PhiReq/phi_stmt_3081/phi_stmt_3081_sources/type_cast_3086/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi24_xx_xcritedgex_xix_xi28_PhiReq/phi_stmt_3081/phi_stmt_3081_sources/type_cast_3086/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi24_xx_xcritedgex_xix_xi28_PhiReq/phi_stmt_3081/phi_stmt_3081_sources/type_cast_3086/SplitProtocol/Sample/rr
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi24_xx_xcritedgex_xix_xi28_PhiReq/phi_stmt_3081/phi_stmt_3081_sources/type_cast_3086/SplitProtocol/Sample/ra
      -- 
    cp_elements(1961) <= cp_elements(1960);
    -- CP-element group 1962 transition  bypass 
    -- predecessors 1960 
    -- successors 1963 
    -- members (4) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi24_xx_xcritedgex_xix_xi28_PhiReq/phi_stmt_3081/phi_stmt_3081_sources/type_cast_3086/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi24_xx_xcritedgex_xix_xi28_PhiReq/phi_stmt_3081/phi_stmt_3081_sources/type_cast_3086/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi24_xx_xcritedgex_xix_xi28_PhiReq/phi_stmt_3081/phi_stmt_3081_sources/type_cast_3086/SplitProtocol/Update/cr
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi24_xx_xcritedgex_xix_xi28_PhiReq/phi_stmt_3081/phi_stmt_3081_sources/type_cast_3086/SplitProtocol/Update/ca
      -- 
    cp_elements(1962) <= cp_elements(1960);
    -- CP-element group 1963 join  transition  bypass 
    -- predecessors 1961 1962 
    -- successors 1964 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi24_xx_xcritedgex_xix_xi28_PhiReq/phi_stmt_3081/phi_stmt_3081_sources/type_cast_3086/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi24_xx_xcritedgex_xix_xi28_PhiReq/phi_stmt_3081/phi_stmt_3081_sources/type_cast_3086/SplitProtocol/$exit
      -- 
    cp_element_group_1963: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1963"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1961) & cp_elements(1962);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1963), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1964 join  transition  output  bypass 
    -- predecessors 1959 1963 
    -- successors 1965 
    -- members (3) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi24_xx_xcritedgex_xix_xi28_PhiReq/phi_stmt_3081/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi24_xx_xcritedgex_xix_xi28_PhiReq/phi_stmt_3081/phi_stmt_3081_sources/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi24_xx_xcritedgex_xix_xi28_PhiReq/phi_stmt_3081/phi_stmt_3081_req
      -- 
    cp_element_group_1964: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1964"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1959) & cp_elements(1963);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1964), clk => clk, reset => reset); --
    end block;
    phi_stmt_3081_req_18184_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1964), ack => phi_stmt_3081_req_0); -- 
    -- CP-element group 1965 join  transition  bypass 
    -- predecessors 1952 1964 
    -- successors 1966 
    -- members (1) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi24_xx_xcritedgex_xix_xi28_PhiReq/$exit
      -- 
    cp_element_group_1965: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1965"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1952) & cp_elements(1964);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1965), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1966 merge  place  bypass 
    -- predecessors 1939 1965 
    -- successors 1967 
    -- members (1) 
      -- 	branch_block_stmt_2042/merge_stmt_3074_PhiReqMerge
      -- 
    cp_elements(1966) <= OrReduce(cp_elements(1939) & cp_elements(1965));
    -- CP-element group 1967 fork  transition  bypass 
    -- predecessors 1966 
    -- successors 1968 1969 
    -- members (1) 
      -- 	branch_block_stmt_2042/merge_stmt_3074_PhiAck/$entry
      -- 
    cp_elements(1967) <= cp_elements(1966);
    -- CP-element group 1968 transition  input  bypass 
    -- predecessors 1967 
    -- successors 1970 
    -- members (1) 
      -- 	branch_block_stmt_2042/merge_stmt_3074_PhiAck/phi_stmt_3075_ack
      -- 
    phi_stmt_3075_ack_18189_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_3075_ack_0, ack => cp_elements(1968)); -- 
    -- CP-element group 1969 transition  input  bypass 
    -- predecessors 1967 
    -- successors 1970 
    -- members (1) 
      -- 	branch_block_stmt_2042/merge_stmt_3074_PhiAck/phi_stmt_3081_ack
      -- 
    phi_stmt_3081_ack_18190_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_3081_ack_0, ack => cp_elements(1969)); -- 
    -- CP-element group 1970 join  transition  bypass 
    -- predecessors 1968 1969 
    -- successors 42 
    -- members (1) 
      -- 	branch_block_stmt_2042/merge_stmt_3074_PhiAck/$exit
      -- 
    cp_element_group_1970: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1970"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1968) & cp_elements(1969);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1970), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1971 transition  bypass 
    -- predecessors 485 
    -- successors 1973 
    -- members (4) 
      -- 	branch_block_stmt_2042/rotor_flux_calcx_xexit_omega_calcx_xexit_PhiReq/phi_stmt_3122/phi_stmt_3122_sources/type_cast_3125/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_2042/rotor_flux_calcx_xexit_omega_calcx_xexit_PhiReq/phi_stmt_3122/phi_stmt_3122_sources/type_cast_3125/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_2042/rotor_flux_calcx_xexit_omega_calcx_xexit_PhiReq/phi_stmt_3122/phi_stmt_3122_sources/type_cast_3125/SplitProtocol/Sample/rr
      -- 	branch_block_stmt_2042/rotor_flux_calcx_xexit_omega_calcx_xexit_PhiReq/phi_stmt_3122/phi_stmt_3122_sources/type_cast_3125/SplitProtocol/Sample/ra
      -- 
    cp_elements(1971) <= cp_elements(485);
    -- CP-element group 1972 transition  bypass 
    -- predecessors 485 
    -- successors 1973 
    -- members (4) 
      -- 	branch_block_stmt_2042/rotor_flux_calcx_xexit_omega_calcx_xexit_PhiReq/phi_stmt_3122/phi_stmt_3122_sources/type_cast_3125/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_2042/rotor_flux_calcx_xexit_omega_calcx_xexit_PhiReq/phi_stmt_3122/phi_stmt_3122_sources/type_cast_3125/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_2042/rotor_flux_calcx_xexit_omega_calcx_xexit_PhiReq/phi_stmt_3122/phi_stmt_3122_sources/type_cast_3125/SplitProtocol/Update/cr
      -- 	branch_block_stmt_2042/rotor_flux_calcx_xexit_omega_calcx_xexit_PhiReq/phi_stmt_3122/phi_stmt_3122_sources/type_cast_3125/SplitProtocol/Update/ca
      -- 
    cp_elements(1972) <= cp_elements(485);
    -- CP-element group 1973 join  transition  output  bypass 
    -- predecessors 1971 1972 
    -- successors 1979 
    -- members (6) 
      -- 	branch_block_stmt_2042/rotor_flux_calcx_xexit_omega_calcx_xexit_PhiReq/$exit
      -- 	branch_block_stmt_2042/rotor_flux_calcx_xexit_omega_calcx_xexit_PhiReq/phi_stmt_3122/$exit
      -- 	branch_block_stmt_2042/rotor_flux_calcx_xexit_omega_calcx_xexit_PhiReq/phi_stmt_3122/phi_stmt_3122_sources/$exit
      -- 	branch_block_stmt_2042/rotor_flux_calcx_xexit_omega_calcx_xexit_PhiReq/phi_stmt_3122/phi_stmt_3122_sources/type_cast_3125/$exit
      -- 	branch_block_stmt_2042/rotor_flux_calcx_xexit_omega_calcx_xexit_PhiReq/phi_stmt_3122/phi_stmt_3122_sources/type_cast_3125/SplitProtocol/$exit
      -- 	branch_block_stmt_2042/rotor_flux_calcx_xexit_omega_calcx_xexit_PhiReq/phi_stmt_3122/phi_stmt_3122_req
      -- 
    cp_element_group_1973: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1973"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1971) & cp_elements(1972);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1973), clk => clk, reset => reset); --
    end block;
    phi_stmt_3122_req_18216_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1973), ack => phi_stmt_3122_req_1); -- 
    -- CP-element group 1974 transition  output  bypass 
    -- predecessors 722 
    -- successors 1975 
    -- members (2) 
      -- 	branch_block_stmt_2042/xx_xcritedgex_xix_xi28_omega_calcx_xexit_PhiReq/phi_stmt_3122/phi_stmt_3122_sources/type_cast_3125/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_2042/xx_xcritedgex_xix_xi28_omega_calcx_xexit_PhiReq/phi_stmt_3122/phi_stmt_3122_sources/type_cast_3125/SplitProtocol/Sample/rr
      -- 
    cp_elements(1974) <= cp_elements(722);
    rr_18235_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1974), ack => type_cast_3125_inst_req_0); -- 
    -- CP-element group 1975 transition  input  bypass 
    -- predecessors 1974 
    -- successors 1978 
    -- members (2) 
      -- 	branch_block_stmt_2042/xx_xcritedgex_xix_xi28_omega_calcx_xexit_PhiReq/phi_stmt_3122/phi_stmt_3122_sources/type_cast_3125/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_2042/xx_xcritedgex_xix_xi28_omega_calcx_xexit_PhiReq/phi_stmt_3122/phi_stmt_3122_sources/type_cast_3125/SplitProtocol/Sample/ra
      -- 
    ra_18236_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3125_inst_ack_0, ack => cp_elements(1975)); -- 
    -- CP-element group 1976 transition  output  bypass 
    -- predecessors 722 
    -- successors 1977 
    -- members (2) 
      -- 	branch_block_stmt_2042/xx_xcritedgex_xix_xi28_omega_calcx_xexit_PhiReq/phi_stmt_3122/phi_stmt_3122_sources/type_cast_3125/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_2042/xx_xcritedgex_xix_xi28_omega_calcx_xexit_PhiReq/phi_stmt_3122/phi_stmt_3122_sources/type_cast_3125/SplitProtocol/Update/cr
      -- 
    cp_elements(1976) <= cp_elements(722);
    cr_18240_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1976), ack => type_cast_3125_inst_req_1); -- 
    -- CP-element group 1977 transition  input  bypass 
    -- predecessors 1976 
    -- successors 1978 
    -- members (2) 
      -- 	branch_block_stmt_2042/xx_xcritedgex_xix_xi28_omega_calcx_xexit_PhiReq/phi_stmt_3122/phi_stmt_3122_sources/type_cast_3125/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_2042/xx_xcritedgex_xix_xi28_omega_calcx_xexit_PhiReq/phi_stmt_3122/phi_stmt_3122_sources/type_cast_3125/SplitProtocol/Update/ca
      -- 
    ca_18241_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3125_inst_ack_1, ack => cp_elements(1977)); -- 
    -- CP-element group 1978 join  transition  output  bypass 
    -- predecessors 1975 1977 
    -- successors 1979 
    -- members (6) 
      -- 	branch_block_stmt_2042/xx_xcritedgex_xix_xi28_omega_calcx_xexit_PhiReq/$exit
      -- 	branch_block_stmt_2042/xx_xcritedgex_xix_xi28_omega_calcx_xexit_PhiReq/phi_stmt_3122/$exit
      -- 	branch_block_stmt_2042/xx_xcritedgex_xix_xi28_omega_calcx_xexit_PhiReq/phi_stmt_3122/phi_stmt_3122_sources/$exit
      -- 	branch_block_stmt_2042/xx_xcritedgex_xix_xi28_omega_calcx_xexit_PhiReq/phi_stmt_3122/phi_stmt_3122_sources/type_cast_3125/$exit
      -- 	branch_block_stmt_2042/xx_xcritedgex_xix_xi28_omega_calcx_xexit_PhiReq/phi_stmt_3122/phi_stmt_3122_sources/type_cast_3125/SplitProtocol/$exit
      -- 	branch_block_stmt_2042/xx_xcritedgex_xix_xi28_omega_calcx_xexit_PhiReq/phi_stmt_3122/phi_stmt_3122_req
      -- 
    cp_element_group_1978: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1978"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1975) & cp_elements(1977);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1978), clk => clk, reset => reset); --
    end block;
    phi_stmt_3122_req_18242_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1978), ack => phi_stmt_3122_req_0); -- 
    -- CP-element group 1979 merge  place  bypass 
    -- predecessors 1973 1978 
    -- successors 1980 
    -- members (1) 
      -- 	branch_block_stmt_2042/merge_stmt_3121_PhiReqMerge
      -- 
    cp_elements(1979) <= OrReduce(cp_elements(1973) & cp_elements(1978));
    -- CP-element group 1980 transition  bypass 
    -- predecessors 1979 
    -- successors 1981 
    -- members (1) 
      -- 	branch_block_stmt_2042/merge_stmt_3121_PhiAck/$entry
      -- 
    cp_elements(1980) <= cp_elements(1979);
    -- CP-element group 1981 transition  place  input  bypass 
    -- predecessors 1980 
    -- successors 723 
    -- members (4) 
      -- 	branch_block_stmt_2042/assign_stmt_3135_to_assign_stmt_3162__entry__
      -- 	branch_block_stmt_2042/merge_stmt_3121__exit__
      -- 	branch_block_stmt_2042/merge_stmt_3121_PhiAck/$exit
      -- 	branch_block_stmt_2042/merge_stmt_3121_PhiAck/phi_stmt_3122_ack
      -- 
    phi_stmt_3122_ack_18247_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_3122_ack_0, ack => cp_elements(1981)); -- 
    -- CP-element group 1982 fork  transition  bypass 
    -- predecessors 46 
    -- successors 1983 1995 
    -- members (1) 
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xix_xix_xpreheader_bbx_xnph7x_xix_xix_xi_PhiReq/$entry
      -- 
    cp_elements(1982) <= cp_elements(46);
    -- CP-element group 1983 fork  transition  bypass 
    -- predecessors 1982 
    -- successors 1984 1988 
    -- members (2) 
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xix_xix_xpreheader_bbx_xnph7x_xix_xix_xi_PhiReq/phi_stmt_3259/$entry
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xix_xix_xpreheader_bbx_xnph7x_xix_xix_xi_PhiReq/phi_stmt_3259/phi_stmt_3259_sources/$entry
      -- 
    cp_elements(1983) <= cp_elements(1982);
    -- CP-element group 1984 fork  transition  bypass 
    -- predecessors 1983 
    -- successors 1985 1986 
    -- members (2) 
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xix_xix_xpreheader_bbx_xnph7x_xix_xix_xi_PhiReq/phi_stmt_3259/phi_stmt_3259_sources/type_cast_3262/$entry
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xix_xix_xpreheader_bbx_xnph7x_xix_xix_xi_PhiReq/phi_stmt_3259/phi_stmt_3259_sources/type_cast_3262/SplitProtocol/$entry
      -- 
    cp_elements(1984) <= cp_elements(1983);
    -- CP-element group 1985 transition  bypass 
    -- predecessors 1984 
    -- successors 1987 
    -- members (4) 
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xix_xix_xpreheader_bbx_xnph7x_xix_xix_xi_PhiReq/phi_stmt_3259/phi_stmt_3259_sources/type_cast_3262/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xix_xix_xpreheader_bbx_xnph7x_xix_xix_xi_PhiReq/phi_stmt_3259/phi_stmt_3259_sources/type_cast_3262/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xix_xix_xpreheader_bbx_xnph7x_xix_xix_xi_PhiReq/phi_stmt_3259/phi_stmt_3259_sources/type_cast_3262/SplitProtocol/Sample/rr
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xix_xix_xpreheader_bbx_xnph7x_xix_xix_xi_PhiReq/phi_stmt_3259/phi_stmt_3259_sources/type_cast_3262/SplitProtocol/Sample/ra
      -- 
    cp_elements(1985) <= cp_elements(1984);
    -- CP-element group 1986 transition  bypass 
    -- predecessors 1984 
    -- successors 1987 
    -- members (4) 
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xix_xix_xpreheader_bbx_xnph7x_xix_xix_xi_PhiReq/phi_stmt_3259/phi_stmt_3259_sources/type_cast_3262/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xix_xix_xpreheader_bbx_xnph7x_xix_xix_xi_PhiReq/phi_stmt_3259/phi_stmt_3259_sources/type_cast_3262/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xix_xix_xpreheader_bbx_xnph7x_xix_xix_xi_PhiReq/phi_stmt_3259/phi_stmt_3259_sources/type_cast_3262/SplitProtocol/Update/cr
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xix_xix_xpreheader_bbx_xnph7x_xix_xix_xi_PhiReq/phi_stmt_3259/phi_stmt_3259_sources/type_cast_3262/SplitProtocol/Update/ca
      -- 
    cp_elements(1986) <= cp_elements(1984);
    -- CP-element group 1987 join  transition  bypass 
    -- predecessors 1985 1986 
    -- successors 1994 
    -- members (2) 
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xix_xix_xpreheader_bbx_xnph7x_xix_xix_xi_PhiReq/phi_stmt_3259/phi_stmt_3259_sources/type_cast_3262/$exit
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xix_xix_xpreheader_bbx_xnph7x_xix_xix_xi_PhiReq/phi_stmt_3259/phi_stmt_3259_sources/type_cast_3262/SplitProtocol/$exit
      -- 
    cp_element_group_1987: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1987"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1985) & cp_elements(1986);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1987), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1988 fork  transition  bypass 
    -- predecessors 1983 
    -- successors 1989 1991 
    -- members (2) 
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xix_xix_xpreheader_bbx_xnph7x_xix_xix_xi_PhiReq/phi_stmt_3259/phi_stmt_3259_sources/type_cast_3264/$entry
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xix_xix_xpreheader_bbx_xnph7x_xix_xix_xi_PhiReq/phi_stmt_3259/phi_stmt_3259_sources/type_cast_3264/SplitProtocol/$entry
      -- 
    cp_elements(1988) <= cp_elements(1983);
    -- CP-element group 1989 transition  output  bypass 
    -- predecessors 1988 
    -- successors 1990 
    -- members (2) 
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xix_xix_xpreheader_bbx_xnph7x_xix_xix_xi_PhiReq/phi_stmt_3259/phi_stmt_3259_sources/type_cast_3264/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xix_xix_xpreheader_bbx_xnph7x_xix_xix_xi_PhiReq/phi_stmt_3259/phi_stmt_3259_sources/type_cast_3264/SplitProtocol/Sample/rr
      -- 
    cp_elements(1989) <= cp_elements(1988);
    rr_18306_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1989), ack => type_cast_3264_inst_req_0); -- 
    -- CP-element group 1990 transition  input  bypass 
    -- predecessors 1989 
    -- successors 1993 
    -- members (2) 
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xix_xix_xpreheader_bbx_xnph7x_xix_xix_xi_PhiReq/phi_stmt_3259/phi_stmt_3259_sources/type_cast_3264/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xix_xix_xpreheader_bbx_xnph7x_xix_xix_xi_PhiReq/phi_stmt_3259/phi_stmt_3259_sources/type_cast_3264/SplitProtocol/Sample/ra
      -- 
    ra_18307_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3264_inst_ack_0, ack => cp_elements(1990)); -- 
    -- CP-element group 1991 transition  output  bypass 
    -- predecessors 1988 
    -- successors 1992 
    -- members (2) 
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xix_xix_xpreheader_bbx_xnph7x_xix_xix_xi_PhiReq/phi_stmt_3259/phi_stmt_3259_sources/type_cast_3264/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xix_xix_xpreheader_bbx_xnph7x_xix_xix_xi_PhiReq/phi_stmt_3259/phi_stmt_3259_sources/type_cast_3264/SplitProtocol/Update/cr
      -- 
    cp_elements(1991) <= cp_elements(1988);
    cr_18311_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1991), ack => type_cast_3264_inst_req_1); -- 
    -- CP-element group 1992 transition  input  bypass 
    -- predecessors 1991 
    -- successors 1993 
    -- members (2) 
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xix_xix_xpreheader_bbx_xnph7x_xix_xix_xi_PhiReq/phi_stmt_3259/phi_stmt_3259_sources/type_cast_3264/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xix_xix_xpreheader_bbx_xnph7x_xix_xix_xi_PhiReq/phi_stmt_3259/phi_stmt_3259_sources/type_cast_3264/SplitProtocol/Update/ca
      -- 
    ca_18312_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3264_inst_ack_1, ack => cp_elements(1992)); -- 
    -- CP-element group 1993 join  transition  bypass 
    -- predecessors 1990 1992 
    -- successors 1994 
    -- members (2) 
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xix_xix_xpreheader_bbx_xnph7x_xix_xix_xi_PhiReq/phi_stmt_3259/phi_stmt_3259_sources/type_cast_3264/$exit
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xix_xix_xpreheader_bbx_xnph7x_xix_xix_xi_PhiReq/phi_stmt_3259/phi_stmt_3259_sources/type_cast_3264/SplitProtocol/$exit
      -- 
    cp_element_group_1993: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1993"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1990) & cp_elements(1992);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1993), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1994 join  transition  output  bypass 
    -- predecessors 1987 1993 
    -- successors 1999 
    -- members (3) 
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xix_xix_xpreheader_bbx_xnph7x_xix_xix_xi_PhiReq/phi_stmt_3259/$exit
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xix_xix_xpreheader_bbx_xnph7x_xix_xix_xi_PhiReq/phi_stmt_3259/phi_stmt_3259_sources/$exit
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xix_xix_xpreheader_bbx_xnph7x_xix_xix_xi_PhiReq/phi_stmt_3259/phi_stmt_3259_req
      -- 
    cp_element_group_1994: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1994"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1987) & cp_elements(1993);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1994), clk => clk, reset => reset); --
    end block;
    phi_stmt_3259_req_18313_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1994), ack => phi_stmt_3259_req_1); -- 
    -- CP-element group 1995 fork  transition  bypass 
    -- predecessors 1982 
    -- successors 1996 1997 
    -- members (4) 
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xix_xix_xpreheader_bbx_xnph7x_xix_xix_xi_PhiReq/phi_stmt_3265/$entry
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xix_xix_xpreheader_bbx_xnph7x_xix_xix_xi_PhiReq/phi_stmt_3265/phi_stmt_3265_sources/$entry
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xix_xix_xpreheader_bbx_xnph7x_xix_xix_xi_PhiReq/phi_stmt_3265/phi_stmt_3265_sources/type_cast_3268/$entry
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xix_xix_xpreheader_bbx_xnph7x_xix_xix_xi_PhiReq/phi_stmt_3265/phi_stmt_3265_sources/type_cast_3268/SplitProtocol/$entry
      -- 
    cp_elements(1995) <= cp_elements(1982);
    -- CP-element group 1996 transition  bypass 
    -- predecessors 1995 
    -- successors 1998 
    -- members (4) 
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xix_xix_xpreheader_bbx_xnph7x_xix_xix_xi_PhiReq/phi_stmt_3265/phi_stmt_3265_sources/type_cast_3268/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xix_xix_xpreheader_bbx_xnph7x_xix_xix_xi_PhiReq/phi_stmt_3265/phi_stmt_3265_sources/type_cast_3268/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xix_xix_xpreheader_bbx_xnph7x_xix_xix_xi_PhiReq/phi_stmt_3265/phi_stmt_3265_sources/type_cast_3268/SplitProtocol/Sample/rr
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xix_xix_xpreheader_bbx_xnph7x_xix_xix_xi_PhiReq/phi_stmt_3265/phi_stmt_3265_sources/type_cast_3268/SplitProtocol/Sample/ra
      -- 
    cp_elements(1996) <= cp_elements(1995);
    -- CP-element group 1997 transition  bypass 
    -- predecessors 1995 
    -- successors 1998 
    -- members (4) 
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xix_xix_xpreheader_bbx_xnph7x_xix_xix_xi_PhiReq/phi_stmt_3265/phi_stmt_3265_sources/type_cast_3268/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xix_xix_xpreheader_bbx_xnph7x_xix_xix_xi_PhiReq/phi_stmt_3265/phi_stmt_3265_sources/type_cast_3268/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xix_xix_xpreheader_bbx_xnph7x_xix_xix_xi_PhiReq/phi_stmt_3265/phi_stmt_3265_sources/type_cast_3268/SplitProtocol/Update/cr
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xix_xix_xpreheader_bbx_xnph7x_xix_xix_xi_PhiReq/phi_stmt_3265/phi_stmt_3265_sources/type_cast_3268/SplitProtocol/Update/ca
      -- 
    cp_elements(1997) <= cp_elements(1995);
    -- CP-element group 1998 join  transition  output  bypass 
    -- predecessors 1996 1997 
    -- successors 1999 
    -- members (5) 
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xix_xix_xpreheader_bbx_xnph7x_xix_xix_xi_PhiReq/phi_stmt_3265/$exit
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xix_xix_xpreheader_bbx_xnph7x_xix_xix_xi_PhiReq/phi_stmt_3265/phi_stmt_3265_sources/$exit
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xix_xix_xpreheader_bbx_xnph7x_xix_xix_xi_PhiReq/phi_stmt_3265/phi_stmt_3265_sources/type_cast_3268/$exit
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xix_xix_xpreheader_bbx_xnph7x_xix_xix_xi_PhiReq/phi_stmt_3265/phi_stmt_3265_sources/type_cast_3268/SplitProtocol/$exit
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xix_xix_xpreheader_bbx_xnph7x_xix_xix_xi_PhiReq/phi_stmt_3265/phi_stmt_3265_req
      -- 
    cp_element_group_1998: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1998"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1996) & cp_elements(1997);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1998), clk => clk, reset => reset); --
    end block;
    phi_stmt_3265_req_18336_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1998), ack => phi_stmt_3265_req_1); -- 
    -- CP-element group 1999 join  transition  bypass 
    -- predecessors 1994 1998 
    -- successors 2020 
    -- members (1) 
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xix_xix_xpreheader_bbx_xnph7x_xix_xix_xi_PhiReq/$exit
      -- 
    cp_element_group_1999: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1999"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1994) & cp_elements(1998);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1999), clk => clk, reset => reset); --
    end block;
    -- CP-element group 2000 fork  transition  bypass 
    -- predecessors 891 
    -- successors 2001 2013 
    -- members (1) 
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi_bbx_xnph7x_xix_xix_xi_PhiReq/$entry
      -- 
    cp_elements(2000) <= cp_elements(891);
    -- CP-element group 2001 fork  transition  bypass 
    -- predecessors 2000 
    -- successors 2002 2008 
    -- members (2) 
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi_bbx_xnph7x_xix_xix_xi_PhiReq/phi_stmt_3259/$entry
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi_bbx_xnph7x_xix_xix_xi_PhiReq/phi_stmt_3259/phi_stmt_3259_sources/$entry
      -- 
    cp_elements(2001) <= cp_elements(2000);
    -- CP-element group 2002 fork  transition  bypass 
    -- predecessors 2001 
    -- successors 2003 2005 
    -- members (2) 
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi_bbx_xnph7x_xix_xix_xi_PhiReq/phi_stmt_3259/phi_stmt_3259_sources/type_cast_3262/$entry
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi_bbx_xnph7x_xix_xix_xi_PhiReq/phi_stmt_3259/phi_stmt_3259_sources/type_cast_3262/SplitProtocol/$entry
      -- 
    cp_elements(2002) <= cp_elements(2001);
    -- CP-element group 2003 transition  output  bypass 
    -- predecessors 2002 
    -- successors 2004 
    -- members (2) 
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi_bbx_xnph7x_xix_xix_xi_PhiReq/phi_stmt_3259/phi_stmt_3259_sources/type_cast_3262/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi_bbx_xnph7x_xix_xix_xi_PhiReq/phi_stmt_3259/phi_stmt_3259_sources/type_cast_3262/SplitProtocol/Sample/rr
      -- 
    cp_elements(2003) <= cp_elements(2002);
    rr_18355_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2003), ack => type_cast_3262_inst_req_0); -- 
    -- CP-element group 2004 transition  input  bypass 
    -- predecessors 2003 
    -- successors 2007 
    -- members (2) 
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi_bbx_xnph7x_xix_xix_xi_PhiReq/phi_stmt_3259/phi_stmt_3259_sources/type_cast_3262/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi_bbx_xnph7x_xix_xix_xi_PhiReq/phi_stmt_3259/phi_stmt_3259_sources/type_cast_3262/SplitProtocol/Sample/ra
      -- 
    ra_18356_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3262_inst_ack_0, ack => cp_elements(2004)); -- 
    -- CP-element group 2005 transition  output  bypass 
    -- predecessors 2002 
    -- successors 2006 
    -- members (2) 
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi_bbx_xnph7x_xix_xix_xi_PhiReq/phi_stmt_3259/phi_stmt_3259_sources/type_cast_3262/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi_bbx_xnph7x_xix_xix_xi_PhiReq/phi_stmt_3259/phi_stmt_3259_sources/type_cast_3262/SplitProtocol/Update/cr
      -- 
    cp_elements(2005) <= cp_elements(2002);
    cr_18360_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2005), ack => type_cast_3262_inst_req_1); -- 
    -- CP-element group 2006 transition  input  bypass 
    -- predecessors 2005 
    -- successors 2007 
    -- members (2) 
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi_bbx_xnph7x_xix_xix_xi_PhiReq/phi_stmt_3259/phi_stmt_3259_sources/type_cast_3262/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi_bbx_xnph7x_xix_xix_xi_PhiReq/phi_stmt_3259/phi_stmt_3259_sources/type_cast_3262/SplitProtocol/Update/ca
      -- 
    ca_18361_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3262_inst_ack_1, ack => cp_elements(2006)); -- 
    -- CP-element group 2007 join  transition  bypass 
    -- predecessors 2004 2006 
    -- successors 2012 
    -- members (2) 
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi_bbx_xnph7x_xix_xix_xi_PhiReq/phi_stmt_3259/phi_stmt_3259_sources/type_cast_3262/$exit
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi_bbx_xnph7x_xix_xix_xi_PhiReq/phi_stmt_3259/phi_stmt_3259_sources/type_cast_3262/SplitProtocol/$exit
      -- 
    cp_element_group_2007: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_2007"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(2004) & cp_elements(2006);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(2007), clk => clk, reset => reset); --
    end block;
    -- CP-element group 2008 fork  transition  bypass 
    -- predecessors 2001 
    -- successors 2009 2010 
    -- members (2) 
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi_bbx_xnph7x_xix_xix_xi_PhiReq/phi_stmt_3259/phi_stmt_3259_sources/type_cast_3264/$entry
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi_bbx_xnph7x_xix_xix_xi_PhiReq/phi_stmt_3259/phi_stmt_3259_sources/type_cast_3264/SplitProtocol/$entry
      -- 
    cp_elements(2008) <= cp_elements(2001);
    -- CP-element group 2009 transition  bypass 
    -- predecessors 2008 
    -- successors 2011 
    -- members (4) 
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi_bbx_xnph7x_xix_xix_xi_PhiReq/phi_stmt_3259/phi_stmt_3259_sources/type_cast_3264/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi_bbx_xnph7x_xix_xix_xi_PhiReq/phi_stmt_3259/phi_stmt_3259_sources/type_cast_3264/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi_bbx_xnph7x_xix_xix_xi_PhiReq/phi_stmt_3259/phi_stmt_3259_sources/type_cast_3264/SplitProtocol/Sample/rr
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi_bbx_xnph7x_xix_xix_xi_PhiReq/phi_stmt_3259/phi_stmt_3259_sources/type_cast_3264/SplitProtocol/Sample/ra
      -- 
    cp_elements(2009) <= cp_elements(2008);
    -- CP-element group 2010 transition  bypass 
    -- predecessors 2008 
    -- successors 2011 
    -- members (4) 
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi_bbx_xnph7x_xix_xix_xi_PhiReq/phi_stmt_3259/phi_stmt_3259_sources/type_cast_3264/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi_bbx_xnph7x_xix_xix_xi_PhiReq/phi_stmt_3259/phi_stmt_3259_sources/type_cast_3264/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi_bbx_xnph7x_xix_xix_xi_PhiReq/phi_stmt_3259/phi_stmt_3259_sources/type_cast_3264/SplitProtocol/Update/cr
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi_bbx_xnph7x_xix_xix_xi_PhiReq/phi_stmt_3259/phi_stmt_3259_sources/type_cast_3264/SplitProtocol/Update/ca
      -- 
    cp_elements(2010) <= cp_elements(2008);
    -- CP-element group 2011 join  transition  bypass 
    -- predecessors 2009 2010 
    -- successors 2012 
    -- members (2) 
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi_bbx_xnph7x_xix_xix_xi_PhiReq/phi_stmt_3259/phi_stmt_3259_sources/type_cast_3264/$exit
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi_bbx_xnph7x_xix_xix_xi_PhiReq/phi_stmt_3259/phi_stmt_3259_sources/type_cast_3264/SplitProtocol/$exit
      -- 
    cp_element_group_2011: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_2011"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(2009) & cp_elements(2010);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(2011), clk => clk, reset => reset); --
    end block;
    -- CP-element group 2012 join  transition  output  bypass 
    -- predecessors 2007 2011 
    -- successors 2019 
    -- members (3) 
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi_bbx_xnph7x_xix_xix_xi_PhiReq/phi_stmt_3259/$exit
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi_bbx_xnph7x_xix_xix_xi_PhiReq/phi_stmt_3259/phi_stmt_3259_sources/$exit
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi_bbx_xnph7x_xix_xix_xi_PhiReq/phi_stmt_3259/phi_stmt_3259_req
      -- 
    cp_element_group_2012: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_2012"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(2007) & cp_elements(2011);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(2012), clk => clk, reset => reset); --
    end block;
    phi_stmt_3259_req_18378_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2012), ack => phi_stmt_3259_req_0); -- 
    -- CP-element group 2013 fork  transition  bypass 
    -- predecessors 2000 
    -- successors 2014 2016 
    -- members (4) 
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi_bbx_xnph7x_xix_xix_xi_PhiReq/phi_stmt_3265/$entry
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi_bbx_xnph7x_xix_xix_xi_PhiReq/phi_stmt_3265/phi_stmt_3265_sources/$entry
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi_bbx_xnph7x_xix_xix_xi_PhiReq/phi_stmt_3265/phi_stmt_3265_sources/type_cast_3268/$entry
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi_bbx_xnph7x_xix_xix_xi_PhiReq/phi_stmt_3265/phi_stmt_3265_sources/type_cast_3268/SplitProtocol/$entry
      -- 
    cp_elements(2013) <= cp_elements(2000);
    -- CP-element group 2014 transition  output  bypass 
    -- predecessors 2013 
    -- successors 2015 
    -- members (2) 
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi_bbx_xnph7x_xix_xix_xi_PhiReq/phi_stmt_3265/phi_stmt_3265_sources/type_cast_3268/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi_bbx_xnph7x_xix_xix_xi_PhiReq/phi_stmt_3265/phi_stmt_3265_sources/type_cast_3268/SplitProtocol/Sample/rr
      -- 
    cp_elements(2014) <= cp_elements(2013);
    rr_18394_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2014), ack => type_cast_3268_inst_req_0); -- 
    -- CP-element group 2015 transition  input  bypass 
    -- predecessors 2014 
    -- successors 2018 
    -- members (2) 
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi_bbx_xnph7x_xix_xix_xi_PhiReq/phi_stmt_3265/phi_stmt_3265_sources/type_cast_3268/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi_bbx_xnph7x_xix_xix_xi_PhiReq/phi_stmt_3265/phi_stmt_3265_sources/type_cast_3268/SplitProtocol/Sample/ra
      -- 
    ra_18395_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3268_inst_ack_0, ack => cp_elements(2015)); -- 
    -- CP-element group 2016 transition  output  bypass 
    -- predecessors 2013 
    -- successors 2017 
    -- members (2) 
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi_bbx_xnph7x_xix_xix_xi_PhiReq/phi_stmt_3265/phi_stmt_3265_sources/type_cast_3268/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi_bbx_xnph7x_xix_xix_xi_PhiReq/phi_stmt_3265/phi_stmt_3265_sources/type_cast_3268/SplitProtocol/Update/cr
      -- 
    cp_elements(2016) <= cp_elements(2013);
    cr_18399_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2016), ack => type_cast_3268_inst_req_1); -- 
    -- CP-element group 2017 transition  input  bypass 
    -- predecessors 2016 
    -- successors 2018 
    -- members (2) 
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi_bbx_xnph7x_xix_xix_xi_PhiReq/phi_stmt_3265/phi_stmt_3265_sources/type_cast_3268/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi_bbx_xnph7x_xix_xix_xi_PhiReq/phi_stmt_3265/phi_stmt_3265_sources/type_cast_3268/SplitProtocol/Update/ca
      -- 
    ca_18400_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3268_inst_ack_1, ack => cp_elements(2017)); -- 
    -- CP-element group 2018 join  transition  output  bypass 
    -- predecessors 2015 2017 
    -- successors 2019 
    -- members (5) 
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi_bbx_xnph7x_xix_xix_xi_PhiReq/phi_stmt_3265/$exit
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi_bbx_xnph7x_xix_xix_xi_PhiReq/phi_stmt_3265/phi_stmt_3265_sources/$exit
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi_bbx_xnph7x_xix_xix_xi_PhiReq/phi_stmt_3265/phi_stmt_3265_sources/type_cast_3268/$exit
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi_bbx_xnph7x_xix_xix_xi_PhiReq/phi_stmt_3265/phi_stmt_3265_sources/type_cast_3268/SplitProtocol/$exit
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi_bbx_xnph7x_xix_xix_xi_PhiReq/phi_stmt_3265/phi_stmt_3265_req
      -- 
    cp_element_group_2018: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_2018"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(2015) & cp_elements(2017);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(2018), clk => clk, reset => reset); --
    end block;
    phi_stmt_3265_req_18401_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2018), ack => phi_stmt_3265_req_0); -- 
    -- CP-element group 2019 join  transition  bypass 
    -- predecessors 2012 2018 
    -- successors 2020 
    -- members (1) 
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi_bbx_xnph7x_xix_xix_xi_PhiReq/$exit
      -- 
    cp_element_group_2019: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_2019"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(2012) & cp_elements(2018);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(2019), clk => clk, reset => reset); --
    end block;
    -- CP-element group 2020 merge  place  bypass 
    -- predecessors 1999 2019 
    -- successors 2021 
    -- members (1) 
      -- 	branch_block_stmt_2042/merge_stmt_3258_PhiReqMerge
      -- 
    cp_elements(2020) <= OrReduce(cp_elements(1999) & cp_elements(2019));
    -- CP-element group 2021 fork  transition  bypass 
    -- predecessors 2020 
    -- successors 2022 2023 
    -- members (1) 
      -- 	branch_block_stmt_2042/merge_stmt_3258_PhiAck/$entry
      -- 
    cp_elements(2021) <= cp_elements(2020);
    -- CP-element group 2022 transition  input  bypass 
    -- predecessors 2021 
    -- successors 2024 
    -- members (1) 
      -- 	branch_block_stmt_2042/merge_stmt_3258_PhiAck/phi_stmt_3259_ack
      -- 
    phi_stmt_3259_ack_18406_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_3259_ack_0, ack => cp_elements(2022)); -- 
    -- CP-element group 2023 transition  input  bypass 
    -- predecessors 2021 
    -- successors 2024 
    -- members (1) 
      -- 	branch_block_stmt_2042/merge_stmt_3258_PhiAck/phi_stmt_3265_ack
      -- 
    phi_stmt_3265_ack_18407_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_3265_ack_0, ack => cp_elements(2023)); -- 
    -- CP-element group 2024 join  transition  bypass 
    -- predecessors 2022 2023 
    -- successors 47 
    -- members (1) 
      -- 	branch_block_stmt_2042/merge_stmt_3258_PhiAck/$exit
      -- 
    cp_element_group_2024: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_2024"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(2022) & cp_elements(2023);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(2024), clk => clk, reset => reset); --
    end block;
    -- CP-element group 2025 fork  transition  bypass 
    -- predecessors 863 
    -- successors 2026 2038 
    -- members (1) 
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi_bbx_xnphx_xix_xix_xi_PhiReq/$entry
      -- 
    cp_elements(2025) <= cp_elements(863);
    -- CP-element group 2026 fork  transition  bypass 
    -- predecessors 2025 
    -- successors 2027 2033 
    -- members (2) 
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi_bbx_xnphx_xix_xix_xi_PhiReq/phi_stmt_3293/$entry
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi_bbx_xnphx_xix_xix_xi_PhiReq/phi_stmt_3293/phi_stmt_3293_sources/$entry
      -- 
    cp_elements(2026) <= cp_elements(2025);
    -- CP-element group 2027 fork  transition  bypass 
    -- predecessors 2026 
    -- successors 2028 2030 
    -- members (2) 
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi_bbx_xnphx_xix_xix_xi_PhiReq/phi_stmt_3293/phi_stmt_3293_sources/type_cast_3296/$entry
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi_bbx_xnphx_xix_xix_xi_PhiReq/phi_stmt_3293/phi_stmt_3293_sources/type_cast_3296/SplitProtocol/$entry
      -- 
    cp_elements(2027) <= cp_elements(2026);
    -- CP-element group 2028 transition  output  bypass 
    -- predecessors 2027 
    -- successors 2029 
    -- members (2) 
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi_bbx_xnphx_xix_xix_xi_PhiReq/phi_stmt_3293/phi_stmt_3293_sources/type_cast_3296/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi_bbx_xnphx_xix_xix_xi_PhiReq/phi_stmt_3293/phi_stmt_3293_sources/type_cast_3296/SplitProtocol/Sample/rr
      -- 
    cp_elements(2028) <= cp_elements(2027);
    rr_18438_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2028), ack => type_cast_3296_inst_req_0); -- 
    -- CP-element group 2029 transition  input  bypass 
    -- predecessors 2028 
    -- successors 2032 
    -- members (2) 
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi_bbx_xnphx_xix_xix_xi_PhiReq/phi_stmt_3293/phi_stmt_3293_sources/type_cast_3296/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi_bbx_xnphx_xix_xix_xi_PhiReq/phi_stmt_3293/phi_stmt_3293_sources/type_cast_3296/SplitProtocol/Sample/ra
      -- 
    ra_18439_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3296_inst_ack_0, ack => cp_elements(2029)); -- 
    -- CP-element group 2030 transition  output  bypass 
    -- predecessors 2027 
    -- successors 2031 
    -- members (2) 
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi_bbx_xnphx_xix_xix_xi_PhiReq/phi_stmt_3293/phi_stmt_3293_sources/type_cast_3296/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi_bbx_xnphx_xix_xix_xi_PhiReq/phi_stmt_3293/phi_stmt_3293_sources/type_cast_3296/SplitProtocol/Update/cr
      -- 
    cp_elements(2030) <= cp_elements(2027);
    cr_18443_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2030), ack => type_cast_3296_inst_req_1); -- 
    -- CP-element group 2031 transition  input  bypass 
    -- predecessors 2030 
    -- successors 2032 
    -- members (2) 
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi_bbx_xnphx_xix_xix_xi_PhiReq/phi_stmt_3293/phi_stmt_3293_sources/type_cast_3296/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi_bbx_xnphx_xix_xix_xi_PhiReq/phi_stmt_3293/phi_stmt_3293_sources/type_cast_3296/SplitProtocol/Update/ca
      -- 
    ca_18444_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3296_inst_ack_1, ack => cp_elements(2031)); -- 
    -- CP-element group 2032 join  transition  bypass 
    -- predecessors 2029 2031 
    -- successors 2037 
    -- members (2) 
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi_bbx_xnphx_xix_xix_xi_PhiReq/phi_stmt_3293/phi_stmt_3293_sources/type_cast_3296/$exit
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi_bbx_xnphx_xix_xix_xi_PhiReq/phi_stmt_3293/phi_stmt_3293_sources/type_cast_3296/SplitProtocol/$exit
      -- 
    cp_element_group_2032: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_2032"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(2029) & cp_elements(2031);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(2032), clk => clk, reset => reset); --
    end block;
    -- CP-element group 2033 fork  transition  bypass 
    -- predecessors 2026 
    -- successors 2034 2035 
    -- members (2) 
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi_bbx_xnphx_xix_xix_xi_PhiReq/phi_stmt_3293/phi_stmt_3293_sources/type_cast_3298/$entry
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi_bbx_xnphx_xix_xix_xi_PhiReq/phi_stmt_3293/phi_stmt_3293_sources/type_cast_3298/SplitProtocol/$entry
      -- 
    cp_elements(2033) <= cp_elements(2026);
    -- CP-element group 2034 transition  bypass 
    -- predecessors 2033 
    -- successors 2036 
    -- members (4) 
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi_bbx_xnphx_xix_xix_xi_PhiReq/phi_stmt_3293/phi_stmt_3293_sources/type_cast_3298/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi_bbx_xnphx_xix_xix_xi_PhiReq/phi_stmt_3293/phi_stmt_3293_sources/type_cast_3298/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi_bbx_xnphx_xix_xix_xi_PhiReq/phi_stmt_3293/phi_stmt_3293_sources/type_cast_3298/SplitProtocol/Sample/rr
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi_bbx_xnphx_xix_xix_xi_PhiReq/phi_stmt_3293/phi_stmt_3293_sources/type_cast_3298/SplitProtocol/Sample/ra
      -- 
    cp_elements(2034) <= cp_elements(2033);
    -- CP-element group 2035 transition  bypass 
    -- predecessors 2033 
    -- successors 2036 
    -- members (4) 
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi_bbx_xnphx_xix_xix_xi_PhiReq/phi_stmt_3293/phi_stmt_3293_sources/type_cast_3298/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi_bbx_xnphx_xix_xix_xi_PhiReq/phi_stmt_3293/phi_stmt_3293_sources/type_cast_3298/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi_bbx_xnphx_xix_xix_xi_PhiReq/phi_stmt_3293/phi_stmt_3293_sources/type_cast_3298/SplitProtocol/Update/cr
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi_bbx_xnphx_xix_xix_xi_PhiReq/phi_stmt_3293/phi_stmt_3293_sources/type_cast_3298/SplitProtocol/Update/ca
      -- 
    cp_elements(2035) <= cp_elements(2033);
    -- CP-element group 2036 join  transition  bypass 
    -- predecessors 2034 2035 
    -- successors 2037 
    -- members (2) 
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi_bbx_xnphx_xix_xix_xi_PhiReq/phi_stmt_3293/phi_stmt_3293_sources/type_cast_3298/$exit
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi_bbx_xnphx_xix_xix_xi_PhiReq/phi_stmt_3293/phi_stmt_3293_sources/type_cast_3298/SplitProtocol/$exit
      -- 
    cp_element_group_2036: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_2036"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(2034) & cp_elements(2035);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(2036), clk => clk, reset => reset); --
    end block;
    -- CP-element group 2037 join  transition  output  bypass 
    -- predecessors 2032 2036 
    -- successors 2044 
    -- members (3) 
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi_bbx_xnphx_xix_xix_xi_PhiReq/phi_stmt_3293/$exit
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi_bbx_xnphx_xix_xix_xi_PhiReq/phi_stmt_3293/phi_stmt_3293_sources/$exit
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi_bbx_xnphx_xix_xix_xi_PhiReq/phi_stmt_3293/phi_stmt_3293_req
      -- 
    cp_element_group_2037: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_2037"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(2032) & cp_elements(2036);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(2037), clk => clk, reset => reset); --
    end block;
    phi_stmt_3293_req_18461_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2037), ack => phi_stmt_3293_req_0); -- 
    -- CP-element group 2038 fork  transition  bypass 
    -- predecessors 2025 
    -- successors 2039 2041 
    -- members (4) 
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi_bbx_xnphx_xix_xix_xi_PhiReq/phi_stmt_3299/$entry
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi_bbx_xnphx_xix_xix_xi_PhiReq/phi_stmt_3299/phi_stmt_3299_sources/$entry
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi_bbx_xnphx_xix_xix_xi_PhiReq/phi_stmt_3299/phi_stmt_3299_sources/type_cast_3302/$entry
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi_bbx_xnphx_xix_xix_xi_PhiReq/phi_stmt_3299/phi_stmt_3299_sources/type_cast_3302/SplitProtocol/$entry
      -- 
    cp_elements(2038) <= cp_elements(2025);
    -- CP-element group 2039 transition  output  bypass 
    -- predecessors 2038 
    -- successors 2040 
    -- members (2) 
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi_bbx_xnphx_xix_xix_xi_PhiReq/phi_stmt_3299/phi_stmt_3299_sources/type_cast_3302/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi_bbx_xnphx_xix_xix_xi_PhiReq/phi_stmt_3299/phi_stmt_3299_sources/type_cast_3302/SplitProtocol/Sample/rr
      -- 
    cp_elements(2039) <= cp_elements(2038);
    rr_18477_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2039), ack => type_cast_3302_inst_req_0); -- 
    -- CP-element group 2040 transition  input  bypass 
    -- predecessors 2039 
    -- successors 2043 
    -- members (2) 
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi_bbx_xnphx_xix_xix_xi_PhiReq/phi_stmt_3299/phi_stmt_3299_sources/type_cast_3302/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi_bbx_xnphx_xix_xix_xi_PhiReq/phi_stmt_3299/phi_stmt_3299_sources/type_cast_3302/SplitProtocol/Sample/ra
      -- 
    ra_18478_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3302_inst_ack_0, ack => cp_elements(2040)); -- 
    -- CP-element group 2041 transition  output  bypass 
    -- predecessors 2038 
    -- successors 2042 
    -- members (2) 
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi_bbx_xnphx_xix_xix_xi_PhiReq/phi_stmt_3299/phi_stmt_3299_sources/type_cast_3302/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi_bbx_xnphx_xix_xix_xi_PhiReq/phi_stmt_3299/phi_stmt_3299_sources/type_cast_3302/SplitProtocol/Update/cr
      -- 
    cp_elements(2041) <= cp_elements(2038);
    cr_18482_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2041), ack => type_cast_3302_inst_req_1); -- 
    -- CP-element group 2042 transition  input  bypass 
    -- predecessors 2041 
    -- successors 2043 
    -- members (2) 
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi_bbx_xnphx_xix_xix_xi_PhiReq/phi_stmt_3299/phi_stmt_3299_sources/type_cast_3302/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi_bbx_xnphx_xix_xix_xi_PhiReq/phi_stmt_3299/phi_stmt_3299_sources/type_cast_3302/SplitProtocol/Update/ca
      -- 
    ca_18483_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3302_inst_ack_1, ack => cp_elements(2042)); -- 
    -- CP-element group 2043 join  transition  output  bypass 
    -- predecessors 2040 2042 
    -- successors 2044 
    -- members (5) 
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi_bbx_xnphx_xix_xix_xi_PhiReq/phi_stmt_3299/$exit
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi_bbx_xnphx_xix_xix_xi_PhiReq/phi_stmt_3299/phi_stmt_3299_sources/$exit
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi_bbx_xnphx_xix_xix_xi_PhiReq/phi_stmt_3299/phi_stmt_3299_sources/type_cast_3302/$exit
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi_bbx_xnphx_xix_xix_xi_PhiReq/phi_stmt_3299/phi_stmt_3299_sources/type_cast_3302/SplitProtocol/$exit
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi_bbx_xnphx_xix_xix_xi_PhiReq/phi_stmt_3299/phi_stmt_3299_req
      -- 
    cp_element_group_2043: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_2043"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(2040) & cp_elements(2042);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(2043), clk => clk, reset => reset); --
    end block;
    phi_stmt_3299_req_18484_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2043), ack => phi_stmt_3299_req_0); -- 
    -- CP-element group 2044 join  transition  bypass 
    -- predecessors 2037 2043 
    -- successors 2063 
    -- members (1) 
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi_bbx_xnphx_xix_xix_xi_PhiReq/$exit
      -- 
    cp_element_group_2044: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_2044"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(2037) & cp_elements(2043);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(2044), clk => clk, reset => reset); --
    end block;
    -- CP-element group 2045 fork  transition  bypass 
    -- predecessors 48 
    -- successors 2046 2058 
    -- members (1) 
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xix_xpreheader_bbx_xnphx_xix_xix_xi_PhiReq/$entry
      -- 
    cp_elements(2045) <= cp_elements(48);
    -- CP-element group 2046 fork  transition  bypass 
    -- predecessors 2045 
    -- successors 2047 2051 
    -- members (2) 
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xix_xpreheader_bbx_xnphx_xix_xix_xi_PhiReq/phi_stmt_3293/$entry
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xix_xpreheader_bbx_xnphx_xix_xix_xi_PhiReq/phi_stmt_3293/phi_stmt_3293_sources/$entry
      -- 
    cp_elements(2046) <= cp_elements(2045);
    -- CP-element group 2047 fork  transition  bypass 
    -- predecessors 2046 
    -- successors 2048 2049 
    -- members (2) 
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xix_xpreheader_bbx_xnphx_xix_xix_xi_PhiReq/phi_stmt_3293/phi_stmt_3293_sources/type_cast_3296/$entry
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xix_xpreheader_bbx_xnphx_xix_xix_xi_PhiReq/phi_stmt_3293/phi_stmt_3293_sources/type_cast_3296/SplitProtocol/$entry
      -- 
    cp_elements(2047) <= cp_elements(2046);
    -- CP-element group 2048 transition  bypass 
    -- predecessors 2047 
    -- successors 2050 
    -- members (4) 
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xix_xpreheader_bbx_xnphx_xix_xix_xi_PhiReq/phi_stmt_3293/phi_stmt_3293_sources/type_cast_3296/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xix_xpreheader_bbx_xnphx_xix_xix_xi_PhiReq/phi_stmt_3293/phi_stmt_3293_sources/type_cast_3296/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xix_xpreheader_bbx_xnphx_xix_xix_xi_PhiReq/phi_stmt_3293/phi_stmt_3293_sources/type_cast_3296/SplitProtocol/Sample/rr
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xix_xpreheader_bbx_xnphx_xix_xix_xi_PhiReq/phi_stmt_3293/phi_stmt_3293_sources/type_cast_3296/SplitProtocol/Sample/ra
      -- 
    cp_elements(2048) <= cp_elements(2047);
    -- CP-element group 2049 transition  bypass 
    -- predecessors 2047 
    -- successors 2050 
    -- members (4) 
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xix_xpreheader_bbx_xnphx_xix_xix_xi_PhiReq/phi_stmt_3293/phi_stmt_3293_sources/type_cast_3296/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xix_xpreheader_bbx_xnphx_xix_xix_xi_PhiReq/phi_stmt_3293/phi_stmt_3293_sources/type_cast_3296/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xix_xpreheader_bbx_xnphx_xix_xix_xi_PhiReq/phi_stmt_3293/phi_stmt_3293_sources/type_cast_3296/SplitProtocol/Update/cr
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xix_xpreheader_bbx_xnphx_xix_xix_xi_PhiReq/phi_stmt_3293/phi_stmt_3293_sources/type_cast_3296/SplitProtocol/Update/ca
      -- 
    cp_elements(2049) <= cp_elements(2047);
    -- CP-element group 2050 join  transition  bypass 
    -- predecessors 2048 2049 
    -- successors 2057 
    -- members (2) 
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xix_xpreheader_bbx_xnphx_xix_xix_xi_PhiReq/phi_stmt_3293/phi_stmt_3293_sources/type_cast_3296/$exit
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xix_xpreheader_bbx_xnphx_xix_xix_xi_PhiReq/phi_stmt_3293/phi_stmt_3293_sources/type_cast_3296/SplitProtocol/$exit
      -- 
    cp_element_group_2050: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_2050"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(2048) & cp_elements(2049);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(2050), clk => clk, reset => reset); --
    end block;
    -- CP-element group 2051 fork  transition  bypass 
    -- predecessors 2046 
    -- successors 2052 2054 
    -- members (2) 
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xix_xpreheader_bbx_xnphx_xix_xix_xi_PhiReq/phi_stmt_3293/phi_stmt_3293_sources/type_cast_3298/$entry
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xix_xpreheader_bbx_xnphx_xix_xix_xi_PhiReq/phi_stmt_3293/phi_stmt_3293_sources/type_cast_3298/SplitProtocol/$entry
      -- 
    cp_elements(2051) <= cp_elements(2046);
    -- CP-element group 2052 transition  output  bypass 
    -- predecessors 2051 
    -- successors 2053 
    -- members (2) 
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xix_xpreheader_bbx_xnphx_xix_xix_xi_PhiReq/phi_stmt_3293/phi_stmt_3293_sources/type_cast_3298/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xix_xpreheader_bbx_xnphx_xix_xix_xi_PhiReq/phi_stmt_3293/phi_stmt_3293_sources/type_cast_3298/SplitProtocol/Sample/rr
      -- 
    cp_elements(2052) <= cp_elements(2051);
    rr_18519_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2052), ack => type_cast_3298_inst_req_0); -- 
    -- CP-element group 2053 transition  input  bypass 
    -- predecessors 2052 
    -- successors 2056 
    -- members (2) 
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xix_xpreheader_bbx_xnphx_xix_xix_xi_PhiReq/phi_stmt_3293/phi_stmt_3293_sources/type_cast_3298/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xix_xpreheader_bbx_xnphx_xix_xix_xi_PhiReq/phi_stmt_3293/phi_stmt_3293_sources/type_cast_3298/SplitProtocol/Sample/ra
      -- 
    ra_18520_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3298_inst_ack_0, ack => cp_elements(2053)); -- 
    -- CP-element group 2054 transition  output  bypass 
    -- predecessors 2051 
    -- successors 2055 
    -- members (2) 
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xix_xpreheader_bbx_xnphx_xix_xix_xi_PhiReq/phi_stmt_3293/phi_stmt_3293_sources/type_cast_3298/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xix_xpreheader_bbx_xnphx_xix_xix_xi_PhiReq/phi_stmt_3293/phi_stmt_3293_sources/type_cast_3298/SplitProtocol/Update/cr
      -- 
    cp_elements(2054) <= cp_elements(2051);
    cr_18524_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2054), ack => type_cast_3298_inst_req_1); -- 
    -- CP-element group 2055 transition  input  bypass 
    -- predecessors 2054 
    -- successors 2056 
    -- members (2) 
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xix_xpreheader_bbx_xnphx_xix_xix_xi_PhiReq/phi_stmt_3293/phi_stmt_3293_sources/type_cast_3298/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xix_xpreheader_bbx_xnphx_xix_xix_xi_PhiReq/phi_stmt_3293/phi_stmt_3293_sources/type_cast_3298/SplitProtocol/Update/ca
      -- 
    ca_18525_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3298_inst_ack_1, ack => cp_elements(2055)); -- 
    -- CP-element group 2056 join  transition  bypass 
    -- predecessors 2053 2055 
    -- successors 2057 
    -- members (2) 
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xix_xpreheader_bbx_xnphx_xix_xix_xi_PhiReq/phi_stmt_3293/phi_stmt_3293_sources/type_cast_3298/$exit
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xix_xpreheader_bbx_xnphx_xix_xix_xi_PhiReq/phi_stmt_3293/phi_stmt_3293_sources/type_cast_3298/SplitProtocol/$exit
      -- 
    cp_element_group_2056: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_2056"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(2053) & cp_elements(2055);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(2056), clk => clk, reset => reset); --
    end block;
    -- CP-element group 2057 join  transition  output  bypass 
    -- predecessors 2050 2056 
    -- successors 2062 
    -- members (3) 
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xix_xpreheader_bbx_xnphx_xix_xix_xi_PhiReq/phi_stmt_3293/$exit
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xix_xpreheader_bbx_xnphx_xix_xix_xi_PhiReq/phi_stmt_3293/phi_stmt_3293_sources/$exit
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xix_xpreheader_bbx_xnphx_xix_xix_xi_PhiReq/phi_stmt_3293/phi_stmt_3293_req
      -- 
    cp_element_group_2057: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_2057"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(2050) & cp_elements(2056);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(2057), clk => clk, reset => reset); --
    end block;
    phi_stmt_3293_req_18526_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2057), ack => phi_stmt_3293_req_1); -- 
    -- CP-element group 2058 fork  transition  bypass 
    -- predecessors 2045 
    -- successors 2059 2060 
    -- members (4) 
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xix_xpreheader_bbx_xnphx_xix_xix_xi_PhiReq/phi_stmt_3299/$entry
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xix_xpreheader_bbx_xnphx_xix_xix_xi_PhiReq/phi_stmt_3299/phi_stmt_3299_sources/$entry
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xix_xpreheader_bbx_xnphx_xix_xix_xi_PhiReq/phi_stmt_3299/phi_stmt_3299_sources/type_cast_3302/$entry
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xix_xpreheader_bbx_xnphx_xix_xix_xi_PhiReq/phi_stmt_3299/phi_stmt_3299_sources/type_cast_3302/SplitProtocol/$entry
      -- 
    cp_elements(2058) <= cp_elements(2045);
    -- CP-element group 2059 transition  bypass 
    -- predecessors 2058 
    -- successors 2061 
    -- members (4) 
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xix_xpreheader_bbx_xnphx_xix_xix_xi_PhiReq/phi_stmt_3299/phi_stmt_3299_sources/type_cast_3302/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xix_xpreheader_bbx_xnphx_xix_xix_xi_PhiReq/phi_stmt_3299/phi_stmt_3299_sources/type_cast_3302/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xix_xpreheader_bbx_xnphx_xix_xix_xi_PhiReq/phi_stmt_3299/phi_stmt_3299_sources/type_cast_3302/SplitProtocol/Sample/rr
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xix_xpreheader_bbx_xnphx_xix_xix_xi_PhiReq/phi_stmt_3299/phi_stmt_3299_sources/type_cast_3302/SplitProtocol/Sample/ra
      -- 
    cp_elements(2059) <= cp_elements(2058);
    -- CP-element group 2060 transition  bypass 
    -- predecessors 2058 
    -- successors 2061 
    -- members (4) 
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xix_xpreheader_bbx_xnphx_xix_xix_xi_PhiReq/phi_stmt_3299/phi_stmt_3299_sources/type_cast_3302/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xix_xpreheader_bbx_xnphx_xix_xix_xi_PhiReq/phi_stmt_3299/phi_stmt_3299_sources/type_cast_3302/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xix_xpreheader_bbx_xnphx_xix_xix_xi_PhiReq/phi_stmt_3299/phi_stmt_3299_sources/type_cast_3302/SplitProtocol/Update/cr
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xix_xpreheader_bbx_xnphx_xix_xix_xi_PhiReq/phi_stmt_3299/phi_stmt_3299_sources/type_cast_3302/SplitProtocol/Update/ca
      -- 
    cp_elements(2060) <= cp_elements(2058);
    -- CP-element group 2061 join  transition  output  bypass 
    -- predecessors 2059 2060 
    -- successors 2062 
    -- members (5) 
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xix_xpreheader_bbx_xnphx_xix_xix_xi_PhiReq/phi_stmt_3299/$exit
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xix_xpreheader_bbx_xnphx_xix_xix_xi_PhiReq/phi_stmt_3299/phi_stmt_3299_sources/$exit
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xix_xpreheader_bbx_xnphx_xix_xix_xi_PhiReq/phi_stmt_3299/phi_stmt_3299_sources/type_cast_3302/$exit
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xix_xpreheader_bbx_xnphx_xix_xix_xi_PhiReq/phi_stmt_3299/phi_stmt_3299_sources/type_cast_3302/SplitProtocol/$exit
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xix_xpreheader_bbx_xnphx_xix_xix_xi_PhiReq/phi_stmt_3299/phi_stmt_3299_req
      -- 
    cp_element_group_2061: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_2061"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(2059) & cp_elements(2060);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(2061), clk => clk, reset => reset); --
    end block;
    phi_stmt_3299_req_18549_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2061), ack => phi_stmt_3299_req_1); -- 
    -- CP-element group 2062 join  transition  bypass 
    -- predecessors 2057 2061 
    -- successors 2063 
    -- members (1) 
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xix_xpreheader_bbx_xnphx_xix_xix_xi_PhiReq/$exit
      -- 
    cp_element_group_2062: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_2062"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(2057) & cp_elements(2061);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(2062), clk => clk, reset => reset); --
    end block;
    -- CP-element group 2063 merge  place  bypass 
    -- predecessors 2044 2062 
    -- successors 2064 
    -- members (1) 
      -- 	branch_block_stmt_2042/merge_stmt_3292_PhiReqMerge
      -- 
    cp_elements(2063) <= OrReduce(cp_elements(2044) & cp_elements(2062));
    -- CP-element group 2064 fork  transition  bypass 
    -- predecessors 2063 
    -- successors 2065 2066 
    -- members (1) 
      -- 	branch_block_stmt_2042/merge_stmt_3292_PhiAck/$entry
      -- 
    cp_elements(2064) <= cp_elements(2063);
    -- CP-element group 2065 transition  input  bypass 
    -- predecessors 2064 
    -- successors 2067 
    -- members (1) 
      -- 	branch_block_stmt_2042/merge_stmt_3292_PhiAck/phi_stmt_3293_ack
      -- 
    phi_stmt_3293_ack_18554_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_3293_ack_0, ack => cp_elements(2065)); -- 
    -- CP-element group 2066 transition  input  bypass 
    -- predecessors 2064 
    -- successors 2067 
    -- members (1) 
      -- 	branch_block_stmt_2042/merge_stmt_3292_PhiAck/phi_stmt_3299_ack
      -- 
    phi_stmt_3299_ack_18555_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_3299_ack_0, ack => cp_elements(2066)); -- 
    -- CP-element group 2067 join  transition  bypass 
    -- predecessors 2065 2066 
    -- successors 49 
    -- members (1) 
      -- 	branch_block_stmt_2042/merge_stmt_3292_PhiAck/$exit
      -- 
    cp_element_group_2067: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_2067"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(2065) & cp_elements(2066);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(2067), clk => clk, reset => reset); --
    end block;
    -- CP-element group 2068 fork  transition  bypass 
    -- predecessors 865 
    -- successors 2069 2075 
    -- members (1) 
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi_xx_x_crit_edgex_xix_xix_xix_xloopexit_PhiReq/$entry
      -- 
    cp_elements(2068) <= cp_elements(865);
    -- CP-element group 2069 fork  transition  bypass 
    -- predecessors 2068 
    -- successors 2070 2072 
    -- members (4) 
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi_xx_x_crit_edgex_xix_xix_xix_xloopexit_PhiReq/phi_stmt_3335/$entry
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi_xx_x_crit_edgex_xix_xix_xix_xloopexit_PhiReq/phi_stmt_3335/phi_stmt_3335_sources/$entry
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi_xx_x_crit_edgex_xix_xix_xix_xloopexit_PhiReq/phi_stmt_3335/phi_stmt_3335_sources/type_cast_3338/$entry
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi_xx_x_crit_edgex_xix_xix_xix_xloopexit_PhiReq/phi_stmt_3335/phi_stmt_3335_sources/type_cast_3338/SplitProtocol/$entry
      -- 
    cp_elements(2069) <= cp_elements(2068);
    -- CP-element group 2070 transition  output  bypass 
    -- predecessors 2069 
    -- successors 2071 
    -- members (2) 
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi_xx_x_crit_edgex_xix_xix_xix_xloopexit_PhiReq/phi_stmt_3335/phi_stmt_3335_sources/type_cast_3338/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi_xx_x_crit_edgex_xix_xix_xix_xloopexit_PhiReq/phi_stmt_3335/phi_stmt_3335_sources/type_cast_3338/SplitProtocol/Sample/rr
      -- 
    cp_elements(2070) <= cp_elements(2069);
    rr_18578_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2070), ack => type_cast_3338_inst_req_0); -- 
    -- CP-element group 2071 transition  input  bypass 
    -- predecessors 2070 
    -- successors 2074 
    -- members (2) 
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi_xx_x_crit_edgex_xix_xix_xix_xloopexit_PhiReq/phi_stmt_3335/phi_stmt_3335_sources/type_cast_3338/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi_xx_x_crit_edgex_xix_xix_xix_xloopexit_PhiReq/phi_stmt_3335/phi_stmt_3335_sources/type_cast_3338/SplitProtocol/Sample/ra
      -- 
    ra_18579_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3338_inst_ack_0, ack => cp_elements(2071)); -- 
    -- CP-element group 2072 transition  output  bypass 
    -- predecessors 2069 
    -- successors 2073 
    -- members (2) 
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi_xx_x_crit_edgex_xix_xix_xix_xloopexit_PhiReq/phi_stmt_3335/phi_stmt_3335_sources/type_cast_3338/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi_xx_x_crit_edgex_xix_xix_xix_xloopexit_PhiReq/phi_stmt_3335/phi_stmt_3335_sources/type_cast_3338/SplitProtocol/Update/cr
      -- 
    cp_elements(2072) <= cp_elements(2069);
    cr_18583_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2072), ack => type_cast_3338_inst_req_1); -- 
    -- CP-element group 2073 transition  input  bypass 
    -- predecessors 2072 
    -- successors 2074 
    -- members (2) 
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi_xx_x_crit_edgex_xix_xix_xix_xloopexit_PhiReq/phi_stmt_3335/phi_stmt_3335_sources/type_cast_3338/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi_xx_x_crit_edgex_xix_xix_xix_xloopexit_PhiReq/phi_stmt_3335/phi_stmt_3335_sources/type_cast_3338/SplitProtocol/Update/ca
      -- 
    ca_18584_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3338_inst_ack_1, ack => cp_elements(2073)); -- 
    -- CP-element group 2074 join  transition  output  bypass 
    -- predecessors 2071 2073 
    -- successors 2081 
    -- members (5) 
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi_xx_x_crit_edgex_xix_xix_xix_xloopexit_PhiReq/phi_stmt_3335/$exit
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi_xx_x_crit_edgex_xix_xix_xix_xloopexit_PhiReq/phi_stmt_3335/phi_stmt_3335_sources/$exit
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi_xx_x_crit_edgex_xix_xix_xix_xloopexit_PhiReq/phi_stmt_3335/phi_stmt_3335_sources/type_cast_3338/$exit
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi_xx_x_crit_edgex_xix_xix_xix_xloopexit_PhiReq/phi_stmt_3335/phi_stmt_3335_sources/type_cast_3338/SplitProtocol/$exit
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi_xx_x_crit_edgex_xix_xix_xix_xloopexit_PhiReq/phi_stmt_3335/phi_stmt_3335_req
      -- 
    cp_element_group_2074: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_2074"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(2071) & cp_elements(2073);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(2074), clk => clk, reset => reset); --
    end block;
    phi_stmt_3335_req_18585_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2074), ack => phi_stmt_3335_req_0); -- 
    -- CP-element group 2075 fork  transition  bypass 
    -- predecessors 2068 
    -- successors 2076 2078 
    -- members (4) 
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi_xx_x_crit_edgex_xix_xix_xix_xloopexit_PhiReq/phi_stmt_3331/$entry
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi_xx_x_crit_edgex_xix_xix_xix_xloopexit_PhiReq/phi_stmt_3331/phi_stmt_3331_sources/$entry
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi_xx_x_crit_edgex_xix_xix_xix_xloopexit_PhiReq/phi_stmt_3331/phi_stmt_3331_sources/type_cast_3334/$entry
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi_xx_x_crit_edgex_xix_xix_xix_xloopexit_PhiReq/phi_stmt_3331/phi_stmt_3331_sources/type_cast_3334/SplitProtocol/$entry
      -- 
    cp_elements(2075) <= cp_elements(2068);
    -- CP-element group 2076 transition  output  bypass 
    -- predecessors 2075 
    -- successors 2077 
    -- members (2) 
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi_xx_x_crit_edgex_xix_xix_xix_xloopexit_PhiReq/phi_stmt_3331/phi_stmt_3331_sources/type_cast_3334/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi_xx_x_crit_edgex_xix_xix_xix_xloopexit_PhiReq/phi_stmt_3331/phi_stmt_3331_sources/type_cast_3334/SplitProtocol/Sample/rr
      -- 
    cp_elements(2076) <= cp_elements(2075);
    rr_18601_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2076), ack => type_cast_3334_inst_req_0); -- 
    -- CP-element group 2077 transition  input  bypass 
    -- predecessors 2076 
    -- successors 2080 
    -- members (2) 
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi_xx_x_crit_edgex_xix_xix_xix_xloopexit_PhiReq/phi_stmt_3331/phi_stmt_3331_sources/type_cast_3334/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi_xx_x_crit_edgex_xix_xix_xix_xloopexit_PhiReq/phi_stmt_3331/phi_stmt_3331_sources/type_cast_3334/SplitProtocol/Sample/ra
      -- 
    ra_18602_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3334_inst_ack_0, ack => cp_elements(2077)); -- 
    -- CP-element group 2078 transition  output  bypass 
    -- predecessors 2075 
    -- successors 2079 
    -- members (2) 
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi_xx_x_crit_edgex_xix_xix_xix_xloopexit_PhiReq/phi_stmt_3331/phi_stmt_3331_sources/type_cast_3334/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi_xx_x_crit_edgex_xix_xix_xix_xloopexit_PhiReq/phi_stmt_3331/phi_stmt_3331_sources/type_cast_3334/SplitProtocol/Update/cr
      -- 
    cp_elements(2078) <= cp_elements(2075);
    cr_18606_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2078), ack => type_cast_3334_inst_req_1); -- 
    -- CP-element group 2079 transition  input  bypass 
    -- predecessors 2078 
    -- successors 2080 
    -- members (2) 
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi_xx_x_crit_edgex_xix_xix_xix_xloopexit_PhiReq/phi_stmt_3331/phi_stmt_3331_sources/type_cast_3334/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi_xx_x_crit_edgex_xix_xix_xix_xloopexit_PhiReq/phi_stmt_3331/phi_stmt_3331_sources/type_cast_3334/SplitProtocol/Update/ca
      -- 
    ca_18607_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3334_inst_ack_1, ack => cp_elements(2079)); -- 
    -- CP-element group 2080 join  transition  output  bypass 
    -- predecessors 2077 2079 
    -- successors 2081 
    -- members (5) 
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi_xx_x_crit_edgex_xix_xix_xix_xloopexit_PhiReq/phi_stmt_3331/$exit
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi_xx_x_crit_edgex_xix_xix_xix_xloopexit_PhiReq/phi_stmt_3331/phi_stmt_3331_sources/$exit
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi_xx_x_crit_edgex_xix_xix_xix_xloopexit_PhiReq/phi_stmt_3331/phi_stmt_3331_sources/type_cast_3334/$exit
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi_xx_x_crit_edgex_xix_xix_xix_xloopexit_PhiReq/phi_stmt_3331/phi_stmt_3331_sources/type_cast_3334/SplitProtocol/$exit
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi_xx_x_crit_edgex_xix_xix_xix_xloopexit_PhiReq/phi_stmt_3331/phi_stmt_3331_req
      -- 
    cp_element_group_2080: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_2080"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(2077) & cp_elements(2079);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(2080), clk => clk, reset => reset); --
    end block;
    phi_stmt_3331_req_18608_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2080), ack => phi_stmt_3331_req_0); -- 
    -- CP-element group 2081 join  transition  bypass 
    -- predecessors 2074 2080 
    -- successors 2082 
    -- members (1) 
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xi_xx_x_crit_edgex_xix_xix_xix_xloopexit_PhiReq/$exit
      -- 
    cp_element_group_2081: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_2081"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(2074) & cp_elements(2080);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(2081), clk => clk, reset => reset); --
    end block;
    -- CP-element group 2082 place  bypass 
    -- predecessors 2081 
    -- successors 2083 
    -- members (1) 
      -- 	branch_block_stmt_2042/merge_stmt_3330_PhiReqMerge
      -- 
    cp_elements(2082) <= cp_elements(2081);
    -- CP-element group 2083 fork  transition  bypass 
    -- predecessors 2082 
    -- successors 2084 2085 
    -- members (1) 
      -- 	branch_block_stmt_2042/merge_stmt_3330_PhiAck/$entry
      -- 
    cp_elements(2083) <= cp_elements(2082);
    -- CP-element group 2084 transition  input  bypass 
    -- predecessors 2083 
    -- successors 2086 
    -- members (1) 
      -- 	branch_block_stmt_2042/merge_stmt_3330_PhiAck/phi_stmt_3331_ack
      -- 
    phi_stmt_3331_ack_18613_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_3331_ack_0, ack => cp_elements(2084)); -- 
    -- CP-element group 2085 transition  input  bypass 
    -- predecessors 2083 
    -- successors 2086 
    -- members (1) 
      -- 	branch_block_stmt_2042/merge_stmt_3330_PhiAck/phi_stmt_3335_ack
      -- 
    phi_stmt_3335_ack_18614_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_3335_ack_0, ack => cp_elements(2085)); -- 
    -- CP-element group 2086 join  transition  bypass 
    -- predecessors 2084 2085 
    -- successors 51 
    -- members (1) 
      -- 	branch_block_stmt_2042/merge_stmt_3330_PhiAck/$exit
      -- 
    cp_element_group_2086: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_2086"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(2084) & cp_elements(2085);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(2086), clk => clk, reset => reset); --
    end block;
    -- CP-element group 2087 fork  transition  bypass 
    -- predecessors 843 
    -- successors 2088 2092 
    -- members (1) 
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xix_xi_xx_x_crit_edgex_xix_xix_xi_PhiReq/$entry
      -- 
    cp_elements(2087) <= cp_elements(843);
    -- CP-element group 2088 fork  transition  bypass 
    -- predecessors 2087 
    -- successors 2089 2090 
    -- members (4) 
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xix_xi_xx_x_crit_edgex_xix_xix_xi_PhiReq/phi_stmt_3348/$entry
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xix_xi_xx_x_crit_edgex_xix_xix_xi_PhiReq/phi_stmt_3348/phi_stmt_3348_sources/$entry
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xix_xi_xx_x_crit_edgex_xix_xix_xi_PhiReq/phi_stmt_3348/phi_stmt_3348_sources/type_cast_3354/$entry
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xix_xi_xx_x_crit_edgex_xix_xix_xi_PhiReq/phi_stmt_3348/phi_stmt_3348_sources/type_cast_3354/SplitProtocol/$entry
      -- 
    cp_elements(2088) <= cp_elements(2087);
    -- CP-element group 2089 transition  bypass 
    -- predecessors 2088 
    -- successors 2091 
    -- members (4) 
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xix_xi_xx_x_crit_edgex_xix_xix_xi_PhiReq/phi_stmt_3348/phi_stmt_3348_sources/type_cast_3354/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xix_xi_xx_x_crit_edgex_xix_xix_xi_PhiReq/phi_stmt_3348/phi_stmt_3348_sources/type_cast_3354/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xix_xi_xx_x_crit_edgex_xix_xix_xi_PhiReq/phi_stmt_3348/phi_stmt_3348_sources/type_cast_3354/SplitProtocol/Sample/rr
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xix_xi_xx_x_crit_edgex_xix_xix_xi_PhiReq/phi_stmt_3348/phi_stmt_3348_sources/type_cast_3354/SplitProtocol/Sample/ra
      -- 
    cp_elements(2089) <= cp_elements(2088);
    -- CP-element group 2090 transition  bypass 
    -- predecessors 2088 
    -- successors 2091 
    -- members (4) 
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xix_xi_xx_x_crit_edgex_xix_xix_xi_PhiReq/phi_stmt_3348/phi_stmt_3348_sources/type_cast_3354/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xix_xi_xx_x_crit_edgex_xix_xix_xi_PhiReq/phi_stmt_3348/phi_stmt_3348_sources/type_cast_3354/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xix_xi_xx_x_crit_edgex_xix_xix_xi_PhiReq/phi_stmt_3348/phi_stmt_3348_sources/type_cast_3354/SplitProtocol/Update/cr
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xix_xi_xx_x_crit_edgex_xix_xix_xi_PhiReq/phi_stmt_3348/phi_stmt_3348_sources/type_cast_3354/SplitProtocol/Update/ca
      -- 
    cp_elements(2090) <= cp_elements(2088);
    -- CP-element group 2091 join  transition  output  bypass 
    -- predecessors 2089 2090 
    -- successors 2104 
    -- members (5) 
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xix_xi_xx_x_crit_edgex_xix_xix_xi_PhiReq/phi_stmt_3348/$exit
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xix_xi_xx_x_crit_edgex_xix_xix_xi_PhiReq/phi_stmt_3348/phi_stmt_3348_sources/$exit
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xix_xi_xx_x_crit_edgex_xix_xix_xi_PhiReq/phi_stmt_3348/phi_stmt_3348_sources/type_cast_3354/$exit
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xix_xi_xx_x_crit_edgex_xix_xix_xi_PhiReq/phi_stmt_3348/phi_stmt_3348_sources/type_cast_3354/SplitProtocol/$exit
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xix_xi_xx_x_crit_edgex_xix_xix_xi_PhiReq/phi_stmt_3348/phi_stmt_3348_req
      -- 
    cp_element_group_2091: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_2091"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(2089) & cp_elements(2090);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(2091), clk => clk, reset => reset); --
    end block;
    phi_stmt_3348_req_18640_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2091), ack => phi_stmt_3348_req_0); -- 
    -- CP-element group 2092 fork  transition  bypass 
    -- predecessors 2087 
    -- successors 2093 2099 
    -- members (2) 
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xix_xi_xx_x_crit_edgex_xix_xix_xi_PhiReq/phi_stmt_3342/$entry
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xix_xi_xx_x_crit_edgex_xix_xix_xi_PhiReq/phi_stmt_3342/phi_stmt_3342_sources/$entry
      -- 
    cp_elements(2092) <= cp_elements(2087);
    -- CP-element group 2093 fork  transition  bypass 
    -- predecessors 2092 
    -- successors 2094 2096 
    -- members (2) 
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xix_xi_xx_x_crit_edgex_xix_xix_xi_PhiReq/phi_stmt_3342/phi_stmt_3342_sources/type_cast_3345/$entry
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xix_xi_xx_x_crit_edgex_xix_xix_xi_PhiReq/phi_stmt_3342/phi_stmt_3342_sources/type_cast_3345/SplitProtocol/$entry
      -- 
    cp_elements(2093) <= cp_elements(2092);
    -- CP-element group 2094 transition  output  bypass 
    -- predecessors 2093 
    -- successors 2095 
    -- members (2) 
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xix_xi_xx_x_crit_edgex_xix_xix_xi_PhiReq/phi_stmt_3342/phi_stmt_3342_sources/type_cast_3345/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xix_xi_xx_x_crit_edgex_xix_xix_xi_PhiReq/phi_stmt_3342/phi_stmt_3342_sources/type_cast_3345/SplitProtocol/Sample/rr
      -- 
    cp_elements(2094) <= cp_elements(2093);
    rr_18656_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2094), ack => type_cast_3345_inst_req_0); -- 
    -- CP-element group 2095 transition  input  bypass 
    -- predecessors 2094 
    -- successors 2098 
    -- members (2) 
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xix_xi_xx_x_crit_edgex_xix_xix_xi_PhiReq/phi_stmt_3342/phi_stmt_3342_sources/type_cast_3345/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xix_xi_xx_x_crit_edgex_xix_xix_xi_PhiReq/phi_stmt_3342/phi_stmt_3342_sources/type_cast_3345/SplitProtocol/Sample/ra
      -- 
    ra_18657_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3345_inst_ack_0, ack => cp_elements(2095)); -- 
    -- CP-element group 2096 transition  output  bypass 
    -- predecessors 2093 
    -- successors 2097 
    -- members (2) 
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xix_xi_xx_x_crit_edgex_xix_xix_xi_PhiReq/phi_stmt_3342/phi_stmt_3342_sources/type_cast_3345/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xix_xi_xx_x_crit_edgex_xix_xix_xi_PhiReq/phi_stmt_3342/phi_stmt_3342_sources/type_cast_3345/SplitProtocol/Update/cr
      -- 
    cp_elements(2096) <= cp_elements(2093);
    cr_18661_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2096), ack => type_cast_3345_inst_req_1); -- 
    -- CP-element group 2097 transition  input  bypass 
    -- predecessors 2096 
    -- successors 2098 
    -- members (2) 
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xix_xi_xx_x_crit_edgex_xix_xix_xi_PhiReq/phi_stmt_3342/phi_stmt_3342_sources/type_cast_3345/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xix_xi_xx_x_crit_edgex_xix_xix_xi_PhiReq/phi_stmt_3342/phi_stmt_3342_sources/type_cast_3345/SplitProtocol/Update/ca
      -- 
    ca_18662_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3345_inst_ack_1, ack => cp_elements(2097)); -- 
    -- CP-element group 2098 join  transition  bypass 
    -- predecessors 2095 2097 
    -- successors 2103 
    -- members (2) 
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xix_xi_xx_x_crit_edgex_xix_xix_xi_PhiReq/phi_stmt_3342/phi_stmt_3342_sources/type_cast_3345/$exit
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xix_xi_xx_x_crit_edgex_xix_xix_xi_PhiReq/phi_stmt_3342/phi_stmt_3342_sources/type_cast_3345/SplitProtocol/$exit
      -- 
    cp_element_group_2098: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_2098"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(2095) & cp_elements(2097);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(2098), clk => clk, reset => reset); --
    end block;
    -- CP-element group 2099 fork  transition  bypass 
    -- predecessors 2092 
    -- successors 2100 2101 
    -- members (2) 
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xix_xi_xx_x_crit_edgex_xix_xix_xi_PhiReq/phi_stmt_3342/phi_stmt_3342_sources/type_cast_3347/$entry
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xix_xi_xx_x_crit_edgex_xix_xix_xi_PhiReq/phi_stmt_3342/phi_stmt_3342_sources/type_cast_3347/SplitProtocol/$entry
      -- 
    cp_elements(2099) <= cp_elements(2092);
    -- CP-element group 2100 transition  bypass 
    -- predecessors 2099 
    -- successors 2102 
    -- members (4) 
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xix_xi_xx_x_crit_edgex_xix_xix_xi_PhiReq/phi_stmt_3342/phi_stmt_3342_sources/type_cast_3347/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xix_xi_xx_x_crit_edgex_xix_xix_xi_PhiReq/phi_stmt_3342/phi_stmt_3342_sources/type_cast_3347/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xix_xi_xx_x_crit_edgex_xix_xix_xi_PhiReq/phi_stmt_3342/phi_stmt_3342_sources/type_cast_3347/SplitProtocol/Sample/rr
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xix_xi_xx_x_crit_edgex_xix_xix_xi_PhiReq/phi_stmt_3342/phi_stmt_3342_sources/type_cast_3347/SplitProtocol/Sample/ra
      -- 
    cp_elements(2100) <= cp_elements(2099);
    -- CP-element group 2101 transition  bypass 
    -- predecessors 2099 
    -- successors 2102 
    -- members (4) 
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xix_xi_xx_x_crit_edgex_xix_xix_xi_PhiReq/phi_stmt_3342/phi_stmt_3342_sources/type_cast_3347/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xix_xi_xx_x_crit_edgex_xix_xix_xi_PhiReq/phi_stmt_3342/phi_stmt_3342_sources/type_cast_3347/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xix_xi_xx_x_crit_edgex_xix_xix_xi_PhiReq/phi_stmt_3342/phi_stmt_3342_sources/type_cast_3347/SplitProtocol/Update/cr
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xix_xi_xx_x_crit_edgex_xix_xix_xi_PhiReq/phi_stmt_3342/phi_stmt_3342_sources/type_cast_3347/SplitProtocol/Update/ca
      -- 
    cp_elements(2101) <= cp_elements(2099);
    -- CP-element group 2102 join  transition  bypass 
    -- predecessors 2100 2101 
    -- successors 2103 
    -- members (2) 
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xix_xi_xx_x_crit_edgex_xix_xix_xi_PhiReq/phi_stmt_3342/phi_stmt_3342_sources/type_cast_3347/$exit
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xix_xi_xx_x_crit_edgex_xix_xix_xi_PhiReq/phi_stmt_3342/phi_stmt_3342_sources/type_cast_3347/SplitProtocol/$exit
      -- 
    cp_element_group_2102: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_2102"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(2100) & cp_elements(2101);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(2102), clk => clk, reset => reset); --
    end block;
    -- CP-element group 2103 join  transition  output  bypass 
    -- predecessors 2098 2102 
    -- successors 2104 
    -- members (3) 
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xix_xi_xx_x_crit_edgex_xix_xix_xi_PhiReq/phi_stmt_3342/$exit
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xix_xi_xx_x_crit_edgex_xix_xix_xi_PhiReq/phi_stmt_3342/phi_stmt_3342_sources/$exit
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xix_xi_xx_x_crit_edgex_xix_xix_xi_PhiReq/phi_stmt_3342/phi_stmt_3342_req
      -- 
    cp_element_group_2103: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_2103"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(2098) & cp_elements(2102);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(2103), clk => clk, reset => reset); --
    end block;
    phi_stmt_3342_req_18679_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2103), ack => phi_stmt_3342_req_0); -- 
    -- CP-element group 2104 join  transition  bypass 
    -- predecessors 2091 2103 
    -- successors 2125 
    -- members (1) 
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xix_xi_xx_x_crit_edgex_xix_xix_xi_PhiReq/$exit
      -- 
    cp_element_group_2104: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_2104"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(2091) & cp_elements(2103);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(2104), clk => clk, reset => reset); --
    end block;
    -- CP-element group 2105 fork  transition  bypass 
    -- predecessors 51 
    -- successors 2106 2112 
    -- members (1) 
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xix_xloopexit_xx_x_crit_edgex_xix_xix_xi_PhiReq/$entry
      -- 
    cp_elements(2105) <= cp_elements(51);
    -- CP-element group 2106 fork  transition  bypass 
    -- predecessors 2105 
    -- successors 2107 2109 
    -- members (4) 
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xix_xloopexit_xx_x_crit_edgex_xix_xix_xi_PhiReq/phi_stmt_3348/$entry
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xix_xloopexit_xx_x_crit_edgex_xix_xix_xi_PhiReq/phi_stmt_3348/phi_stmt_3348_sources/$entry
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xix_xloopexit_xx_x_crit_edgex_xix_xix_xi_PhiReq/phi_stmt_3348/phi_stmt_3348_sources/type_cast_3354/$entry
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xix_xloopexit_xx_x_crit_edgex_xix_xix_xi_PhiReq/phi_stmt_3348/phi_stmt_3348_sources/type_cast_3354/SplitProtocol/$entry
      -- 
    cp_elements(2106) <= cp_elements(2105);
    -- CP-element group 2107 transition  output  bypass 
    -- predecessors 2106 
    -- successors 2108 
    -- members (2) 
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xix_xloopexit_xx_x_crit_edgex_xix_xix_xi_PhiReq/phi_stmt_3348/phi_stmt_3348_sources/type_cast_3354/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xix_xloopexit_xx_x_crit_edgex_xix_xix_xi_PhiReq/phi_stmt_3348/phi_stmt_3348_sources/type_cast_3354/SplitProtocol/Sample/rr
      -- 
    cp_elements(2107) <= cp_elements(2106);
    rr_18698_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2107), ack => type_cast_3354_inst_req_0); -- 
    -- CP-element group 2108 transition  input  bypass 
    -- predecessors 2107 
    -- successors 2111 
    -- members (2) 
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xix_xloopexit_xx_x_crit_edgex_xix_xix_xi_PhiReq/phi_stmt_3348/phi_stmt_3348_sources/type_cast_3354/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xix_xloopexit_xx_x_crit_edgex_xix_xix_xi_PhiReq/phi_stmt_3348/phi_stmt_3348_sources/type_cast_3354/SplitProtocol/Sample/ra
      -- 
    ra_18699_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3354_inst_ack_0, ack => cp_elements(2108)); -- 
    -- CP-element group 2109 transition  output  bypass 
    -- predecessors 2106 
    -- successors 2110 
    -- members (2) 
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xix_xloopexit_xx_x_crit_edgex_xix_xix_xi_PhiReq/phi_stmt_3348/phi_stmt_3348_sources/type_cast_3354/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xix_xloopexit_xx_x_crit_edgex_xix_xix_xi_PhiReq/phi_stmt_3348/phi_stmt_3348_sources/type_cast_3354/SplitProtocol/Update/cr
      -- 
    cp_elements(2109) <= cp_elements(2106);
    cr_18703_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2109), ack => type_cast_3354_inst_req_1); -- 
    -- CP-element group 2110 transition  input  bypass 
    -- predecessors 2109 
    -- successors 2111 
    -- members (2) 
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xix_xloopexit_xx_x_crit_edgex_xix_xix_xi_PhiReq/phi_stmt_3348/phi_stmt_3348_sources/type_cast_3354/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xix_xloopexit_xx_x_crit_edgex_xix_xix_xi_PhiReq/phi_stmt_3348/phi_stmt_3348_sources/type_cast_3354/SplitProtocol/Update/ca
      -- 
    ca_18704_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3354_inst_ack_1, ack => cp_elements(2110)); -- 
    -- CP-element group 2111 join  transition  output  bypass 
    -- predecessors 2108 2110 
    -- successors 2124 
    -- members (5) 
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xix_xloopexit_xx_x_crit_edgex_xix_xix_xi_PhiReq/phi_stmt_3348/$exit
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xix_xloopexit_xx_x_crit_edgex_xix_xix_xi_PhiReq/phi_stmt_3348/phi_stmt_3348_sources/$exit
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xix_xloopexit_xx_x_crit_edgex_xix_xix_xi_PhiReq/phi_stmt_3348/phi_stmt_3348_sources/type_cast_3354/$exit
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xix_xloopexit_xx_x_crit_edgex_xix_xix_xi_PhiReq/phi_stmt_3348/phi_stmt_3348_sources/type_cast_3354/SplitProtocol/$exit
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xix_xloopexit_xx_x_crit_edgex_xix_xix_xi_PhiReq/phi_stmt_3348/phi_stmt_3348_req
      -- 
    cp_element_group_2111: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_2111"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(2108) & cp_elements(2110);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(2111), clk => clk, reset => reset); --
    end block;
    phi_stmt_3348_req_18705_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2111), ack => phi_stmt_3348_req_1); -- 
    -- CP-element group 2112 fork  transition  bypass 
    -- predecessors 2105 
    -- successors 2113 2117 
    -- members (2) 
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xix_xloopexit_xx_x_crit_edgex_xix_xix_xi_PhiReq/phi_stmt_3342/$entry
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xix_xloopexit_xx_x_crit_edgex_xix_xix_xi_PhiReq/phi_stmt_3342/phi_stmt_3342_sources/$entry
      -- 
    cp_elements(2112) <= cp_elements(2105);
    -- CP-element group 2113 fork  transition  bypass 
    -- predecessors 2112 
    -- successors 2114 2115 
    -- members (2) 
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xix_xloopexit_xx_x_crit_edgex_xix_xix_xi_PhiReq/phi_stmt_3342/phi_stmt_3342_sources/type_cast_3345/$entry
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xix_xloopexit_xx_x_crit_edgex_xix_xix_xi_PhiReq/phi_stmt_3342/phi_stmt_3342_sources/type_cast_3345/SplitProtocol/$entry
      -- 
    cp_elements(2113) <= cp_elements(2112);
    -- CP-element group 2114 transition  bypass 
    -- predecessors 2113 
    -- successors 2116 
    -- members (4) 
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xix_xloopexit_xx_x_crit_edgex_xix_xix_xi_PhiReq/phi_stmt_3342/phi_stmt_3342_sources/type_cast_3345/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xix_xloopexit_xx_x_crit_edgex_xix_xix_xi_PhiReq/phi_stmt_3342/phi_stmt_3342_sources/type_cast_3345/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xix_xloopexit_xx_x_crit_edgex_xix_xix_xi_PhiReq/phi_stmt_3342/phi_stmt_3342_sources/type_cast_3345/SplitProtocol/Sample/rr
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xix_xloopexit_xx_x_crit_edgex_xix_xix_xi_PhiReq/phi_stmt_3342/phi_stmt_3342_sources/type_cast_3345/SplitProtocol/Sample/ra
      -- 
    cp_elements(2114) <= cp_elements(2113);
    -- CP-element group 2115 transition  bypass 
    -- predecessors 2113 
    -- successors 2116 
    -- members (4) 
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xix_xloopexit_xx_x_crit_edgex_xix_xix_xi_PhiReq/phi_stmt_3342/phi_stmt_3342_sources/type_cast_3345/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xix_xloopexit_xx_x_crit_edgex_xix_xix_xi_PhiReq/phi_stmt_3342/phi_stmt_3342_sources/type_cast_3345/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xix_xloopexit_xx_x_crit_edgex_xix_xix_xi_PhiReq/phi_stmt_3342/phi_stmt_3342_sources/type_cast_3345/SplitProtocol/Update/cr
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xix_xloopexit_xx_x_crit_edgex_xix_xix_xi_PhiReq/phi_stmt_3342/phi_stmt_3342_sources/type_cast_3345/SplitProtocol/Update/ca
      -- 
    cp_elements(2115) <= cp_elements(2113);
    -- CP-element group 2116 join  transition  bypass 
    -- predecessors 2114 2115 
    -- successors 2123 
    -- members (2) 
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xix_xloopexit_xx_x_crit_edgex_xix_xix_xi_PhiReq/phi_stmt_3342/phi_stmt_3342_sources/type_cast_3345/$exit
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xix_xloopexit_xx_x_crit_edgex_xix_xix_xi_PhiReq/phi_stmt_3342/phi_stmt_3342_sources/type_cast_3345/SplitProtocol/$exit
      -- 
    cp_element_group_2116: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_2116"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(2114) & cp_elements(2115);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(2116), clk => clk, reset => reset); --
    end block;
    -- CP-element group 2117 fork  transition  bypass 
    -- predecessors 2112 
    -- successors 2118 2120 
    -- members (2) 
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xix_xloopexit_xx_x_crit_edgex_xix_xix_xi_PhiReq/phi_stmt_3342/phi_stmt_3342_sources/type_cast_3347/$entry
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xix_xloopexit_xx_x_crit_edgex_xix_xix_xi_PhiReq/phi_stmt_3342/phi_stmt_3342_sources/type_cast_3347/SplitProtocol/$entry
      -- 
    cp_elements(2117) <= cp_elements(2112);
    -- CP-element group 2118 transition  output  bypass 
    -- predecessors 2117 
    -- successors 2119 
    -- members (2) 
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xix_xloopexit_xx_x_crit_edgex_xix_xix_xi_PhiReq/phi_stmt_3342/phi_stmt_3342_sources/type_cast_3347/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xix_xloopexit_xx_x_crit_edgex_xix_xix_xi_PhiReq/phi_stmt_3342/phi_stmt_3342_sources/type_cast_3347/SplitProtocol/Sample/rr
      -- 
    cp_elements(2118) <= cp_elements(2117);
    rr_18737_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2118), ack => type_cast_3347_inst_req_0); -- 
    -- CP-element group 2119 transition  input  bypass 
    -- predecessors 2118 
    -- successors 2122 
    -- members (2) 
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xix_xloopexit_xx_x_crit_edgex_xix_xix_xi_PhiReq/phi_stmt_3342/phi_stmt_3342_sources/type_cast_3347/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xix_xloopexit_xx_x_crit_edgex_xix_xix_xi_PhiReq/phi_stmt_3342/phi_stmt_3342_sources/type_cast_3347/SplitProtocol/Sample/ra
      -- 
    ra_18738_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3347_inst_ack_0, ack => cp_elements(2119)); -- 
    -- CP-element group 2120 transition  output  bypass 
    -- predecessors 2117 
    -- successors 2121 
    -- members (2) 
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xix_xloopexit_xx_x_crit_edgex_xix_xix_xi_PhiReq/phi_stmt_3342/phi_stmt_3342_sources/type_cast_3347/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xix_xloopexit_xx_x_crit_edgex_xix_xix_xi_PhiReq/phi_stmt_3342/phi_stmt_3342_sources/type_cast_3347/SplitProtocol/Update/cr
      -- 
    cp_elements(2120) <= cp_elements(2117);
    cr_18742_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2120), ack => type_cast_3347_inst_req_1); -- 
    -- CP-element group 2121 transition  input  bypass 
    -- predecessors 2120 
    -- successors 2122 
    -- members (2) 
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xix_xloopexit_xx_x_crit_edgex_xix_xix_xi_PhiReq/phi_stmt_3342/phi_stmt_3342_sources/type_cast_3347/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xix_xloopexit_xx_x_crit_edgex_xix_xix_xi_PhiReq/phi_stmt_3342/phi_stmt_3342_sources/type_cast_3347/SplitProtocol/Update/ca
      -- 
    ca_18743_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3347_inst_ack_1, ack => cp_elements(2121)); -- 
    -- CP-element group 2122 join  transition  bypass 
    -- predecessors 2119 2121 
    -- successors 2123 
    -- members (2) 
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xix_xloopexit_xx_x_crit_edgex_xix_xix_xi_PhiReq/phi_stmt_3342/phi_stmt_3342_sources/type_cast_3347/$exit
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xix_xloopexit_xx_x_crit_edgex_xix_xix_xi_PhiReq/phi_stmt_3342/phi_stmt_3342_sources/type_cast_3347/SplitProtocol/$exit
      -- 
    cp_element_group_2122: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_2122"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(2119) & cp_elements(2121);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(2122), clk => clk, reset => reset); --
    end block;
    -- CP-element group 2123 join  transition  output  bypass 
    -- predecessors 2116 2122 
    -- successors 2124 
    -- members (3) 
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xix_xloopexit_xx_x_crit_edgex_xix_xix_xi_PhiReq/phi_stmt_3342/$exit
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xix_xloopexit_xx_x_crit_edgex_xix_xix_xi_PhiReq/phi_stmt_3342/phi_stmt_3342_sources/$exit
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xix_xloopexit_xx_x_crit_edgex_xix_xix_xi_PhiReq/phi_stmt_3342/phi_stmt_3342_req
      -- 
    cp_element_group_2123: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_2123"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(2116) & cp_elements(2122);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(2123), clk => clk, reset => reset); --
    end block;
    phi_stmt_3342_req_18744_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2123), ack => phi_stmt_3342_req_1); -- 
    -- CP-element group 2124 join  transition  bypass 
    -- predecessors 2111 2123 
    -- successors 2125 
    -- members (1) 
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xix_xloopexit_xx_x_crit_edgex_xix_xix_xi_PhiReq/$exit
      -- 
    cp_element_group_2124: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_2124"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(2111) & cp_elements(2123);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(2124), clk => clk, reset => reset); --
    end block;
    -- CP-element group 2125 merge  place  bypass 
    -- predecessors 2104 2124 
    -- successors 2126 
    -- members (1) 
      -- 	branch_block_stmt_2042/merge_stmt_3341_PhiReqMerge
      -- 
    cp_elements(2125) <= OrReduce(cp_elements(2104) & cp_elements(2124));
    -- CP-element group 2126 fork  transition  bypass 
    -- predecessors 2125 
    -- successors 2127 2128 
    -- members (1) 
      -- 	branch_block_stmt_2042/merge_stmt_3341_PhiAck/$entry
      -- 
    cp_elements(2126) <= cp_elements(2125);
    -- CP-element group 2127 transition  input  bypass 
    -- predecessors 2126 
    -- successors 2129 
    -- members (1) 
      -- 	branch_block_stmt_2042/merge_stmt_3341_PhiAck/phi_stmt_3342_ack
      -- 
    phi_stmt_3342_ack_18749_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_3342_ack_0, ack => cp_elements(2127)); -- 
    -- CP-element group 2128 transition  input  bypass 
    -- predecessors 2126 
    -- successors 2129 
    -- members (1) 
      -- 	branch_block_stmt_2042/merge_stmt_3341_PhiAck/phi_stmt_3348_ack
      -- 
    phi_stmt_3348_ack_18750_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_3348_ack_0, ack => cp_elements(2128)); -- 
    -- CP-element group 2129 join  transition  bypass 
    -- predecessors 2127 2128 
    -- successors 52 
    -- members (1) 
      -- 	branch_block_stmt_2042/merge_stmt_3341_PhiAck/$exit
      -- 
    cp_element_group_2129: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_2129"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(2127) & cp_elements(2128);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(2129), clk => clk, reset => reset); --
    end block;
    -- CP-element group 2130 transition  output  bypass 
    -- predecessors 889 
    -- successors 2131 
    -- members (2) 
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi_xx_xloopexitx_xix_xix_xix_xloopexit_PhiReq/phi_stmt_3378/phi_stmt_3378_sources/type_cast_3381/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi_xx_xloopexitx_xix_xix_xix_xloopexit_PhiReq/phi_stmt_3378/phi_stmt_3378_sources/type_cast_3381/SplitProtocol/Sample/rr
      -- 
    cp_elements(2130) <= cp_elements(889);
    rr_18773_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2130), ack => type_cast_3381_inst_req_0); -- 
    -- CP-element group 2131 transition  input  bypass 
    -- predecessors 2130 
    -- successors 2134 
    -- members (2) 
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi_xx_xloopexitx_xix_xix_xix_xloopexit_PhiReq/phi_stmt_3378/phi_stmt_3378_sources/type_cast_3381/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi_xx_xloopexitx_xix_xix_xix_xloopexit_PhiReq/phi_stmt_3378/phi_stmt_3378_sources/type_cast_3381/SplitProtocol/Sample/ra
      -- 
    ra_18774_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3381_inst_ack_0, ack => cp_elements(2131)); -- 
    -- CP-element group 2132 transition  output  bypass 
    -- predecessors 889 
    -- successors 2133 
    -- members (2) 
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi_xx_xloopexitx_xix_xix_xix_xloopexit_PhiReq/phi_stmt_3378/phi_stmt_3378_sources/type_cast_3381/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi_xx_xloopexitx_xix_xix_xix_xloopexit_PhiReq/phi_stmt_3378/phi_stmt_3378_sources/type_cast_3381/SplitProtocol/Update/cr
      -- 
    cp_elements(2132) <= cp_elements(889);
    cr_18778_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2132), ack => type_cast_3381_inst_req_1); -- 
    -- CP-element group 2133 transition  input  bypass 
    -- predecessors 2132 
    -- successors 2134 
    -- members (2) 
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi_xx_xloopexitx_xix_xix_xix_xloopexit_PhiReq/phi_stmt_3378/phi_stmt_3378_sources/type_cast_3381/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi_xx_xloopexitx_xix_xix_xix_xloopexit_PhiReq/phi_stmt_3378/phi_stmt_3378_sources/type_cast_3381/SplitProtocol/Update/ca
      -- 
    ca_18779_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3381_inst_ack_1, ack => cp_elements(2133)); -- 
    -- CP-element group 2134 join  transition  place  output  bypass 
    -- predecessors 2131 2133 
    -- successors 2135 
    -- members (8) 
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi_xx_xloopexitx_xix_xix_xix_xloopexit_PhiReq/$exit
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi_xx_xloopexitx_xix_xix_xix_xloopexit_PhiReq/phi_stmt_3378/$exit
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi_xx_xloopexitx_xix_xix_xix_xloopexit_PhiReq/phi_stmt_3378/phi_stmt_3378_sources/$exit
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi_xx_xloopexitx_xix_xix_xix_xloopexit_PhiReq/phi_stmt_3378/phi_stmt_3378_sources/type_cast_3381/$exit
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi_xx_xloopexitx_xix_xix_xix_xloopexit_PhiReq/phi_stmt_3378/phi_stmt_3378_sources/type_cast_3381/SplitProtocol/$exit
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xi_xx_xloopexitx_xix_xix_xix_xloopexit_PhiReq/phi_stmt_3378/phi_stmt_3378_req
      -- 	branch_block_stmt_2042/merge_stmt_3377_PhiReqMerge
      -- 	branch_block_stmt_2042/merge_stmt_3377_PhiAck/$entry
      -- 
    cp_element_group_2134: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_2134"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(2131) & cp_elements(2133);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(2134), clk => clk, reset => reset); --
    end block;
    phi_stmt_3378_req_18780_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2134), ack => phi_stmt_3378_req_0); -- 
    -- CP-element group 2135 transition  input  bypass 
    -- predecessors 2134 
    -- successors 54 
    -- members (2) 
      -- 	branch_block_stmt_2042/merge_stmt_3377_PhiAck/$exit
      -- 	branch_block_stmt_2042/merge_stmt_3377_PhiAck/phi_stmt_3378_ack
      -- 
    phi_stmt_3378_ack_18785_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_3378_ack_0, ack => cp_elements(2135)); -- 
    -- CP-element group 2136 transition  bypass 
    -- predecessors 822 
    -- successors 2138 
    -- members (4) 
      -- 	branch_block_stmt_2042/bb_41_xx_xloopexitx_xix_xix_xi_PhiReq/phi_stmt_3385/phi_stmt_3385_sources/type_cast_3391/SplitProtocol/Sample/ra
      -- 	branch_block_stmt_2042/bb_41_xx_xloopexitx_xix_xix_xi_PhiReq/phi_stmt_3385/phi_stmt_3385_sources/type_cast_3391/SplitProtocol/Sample/rr
      -- 	branch_block_stmt_2042/bb_41_xx_xloopexitx_xix_xix_xi_PhiReq/phi_stmt_3385/phi_stmt_3385_sources/type_cast_3391/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_2042/bb_41_xx_xloopexitx_xix_xix_xi_PhiReq/phi_stmt_3385/phi_stmt_3385_sources/type_cast_3391/SplitProtocol/Sample/$entry
      -- 
    cp_elements(2136) <= cp_elements(822);
    -- CP-element group 2137 transition  bypass 
    -- predecessors 822 
    -- successors 2138 
    -- members (4) 
      -- 	branch_block_stmt_2042/bb_41_xx_xloopexitx_xix_xix_xi_PhiReq/phi_stmt_3385/phi_stmt_3385_sources/type_cast_3391/SplitProtocol/Update/ca
      -- 	branch_block_stmt_2042/bb_41_xx_xloopexitx_xix_xix_xi_PhiReq/phi_stmt_3385/phi_stmt_3385_sources/type_cast_3391/SplitProtocol/Update/cr
      -- 	branch_block_stmt_2042/bb_41_xx_xloopexitx_xix_xix_xi_PhiReq/phi_stmt_3385/phi_stmt_3385_sources/type_cast_3391/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_2042/bb_41_xx_xloopexitx_xix_xix_xi_PhiReq/phi_stmt_3385/phi_stmt_3385_sources/type_cast_3391/SplitProtocol/Update/$entry
      -- 
    cp_elements(2137) <= cp_elements(822);
    -- CP-element group 2138 join  transition  output  bypass 
    -- predecessors 2136 2137 
    -- successors 2144 
    -- members (6) 
      -- 	branch_block_stmt_2042/bb_41_xx_xloopexitx_xix_xix_xi_PhiReq/phi_stmt_3385/phi_stmt_3385_req
      -- 	branch_block_stmt_2042/bb_41_xx_xloopexitx_xix_xix_xi_PhiReq/$exit
      -- 	branch_block_stmt_2042/bb_41_xx_xloopexitx_xix_xix_xi_PhiReq/phi_stmt_3385/$exit
      -- 	branch_block_stmt_2042/bb_41_xx_xloopexitx_xix_xix_xi_PhiReq/phi_stmt_3385/phi_stmt_3385_sources/$exit
      -- 	branch_block_stmt_2042/bb_41_xx_xloopexitx_xix_xix_xi_PhiReq/phi_stmt_3385/phi_stmt_3385_sources/type_cast_3391/$exit
      -- 	branch_block_stmt_2042/bb_41_xx_xloopexitx_xix_xix_xi_PhiReq/phi_stmt_3385/phi_stmt_3385_sources/type_cast_3391/SplitProtocol/$exit
      -- 
    cp_element_group_2138: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_2138"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(2136) & cp_elements(2137);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(2138), clk => clk, reset => reset); --
    end block;
    phi_stmt_3385_req_18811_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2138), ack => phi_stmt_3385_req_0); -- 
    -- CP-element group 2139 transition  output  bypass 
    -- predecessors 54 
    -- successors 2140 
    -- members (2) 
      -- 	branch_block_stmt_2042/xx_xloopexitx_xix_xix_xix_xloopexit_xx_xloopexitx_xix_xix_xi_PhiReq/phi_stmt_3385/phi_stmt_3385_sources/type_cast_3391/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_2042/xx_xloopexitx_xix_xix_xix_xloopexit_xx_xloopexitx_xix_xix_xi_PhiReq/phi_stmt_3385/phi_stmt_3385_sources/type_cast_3391/SplitProtocol/Sample/rr
      -- 
    cp_elements(2139) <= cp_elements(54);
    rr_18830_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2139), ack => type_cast_3391_inst_req_0); -- 
    -- CP-element group 2140 transition  input  bypass 
    -- predecessors 2139 
    -- successors 2143 
    -- members (2) 
      -- 	branch_block_stmt_2042/xx_xloopexitx_xix_xix_xix_xloopexit_xx_xloopexitx_xix_xix_xi_PhiReq/phi_stmt_3385/phi_stmt_3385_sources/type_cast_3391/SplitProtocol/Sample/ra
      -- 	branch_block_stmt_2042/xx_xloopexitx_xix_xix_xix_xloopexit_xx_xloopexitx_xix_xix_xi_PhiReq/phi_stmt_3385/phi_stmt_3385_sources/type_cast_3391/SplitProtocol/Sample/$exit
      -- 
    ra_18831_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3391_inst_ack_0, ack => cp_elements(2140)); -- 
    -- CP-element group 2141 transition  output  bypass 
    -- predecessors 54 
    -- successors 2142 
    -- members (2) 
      -- 	branch_block_stmt_2042/xx_xloopexitx_xix_xix_xix_xloopexit_xx_xloopexitx_xix_xix_xi_PhiReq/phi_stmt_3385/phi_stmt_3385_sources/type_cast_3391/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_2042/xx_xloopexitx_xix_xix_xix_xloopexit_xx_xloopexitx_xix_xix_xi_PhiReq/phi_stmt_3385/phi_stmt_3385_sources/type_cast_3391/SplitProtocol/Update/cr
      -- 
    cp_elements(2141) <= cp_elements(54);
    cr_18835_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2141), ack => type_cast_3391_inst_req_1); -- 
    -- CP-element group 2142 transition  input  bypass 
    -- predecessors 2141 
    -- successors 2143 
    -- members (2) 
      -- 	branch_block_stmt_2042/xx_xloopexitx_xix_xix_xix_xloopexit_xx_xloopexitx_xix_xix_xi_PhiReq/phi_stmt_3385/phi_stmt_3385_sources/type_cast_3391/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_2042/xx_xloopexitx_xix_xix_xix_xloopexit_xx_xloopexitx_xix_xix_xi_PhiReq/phi_stmt_3385/phi_stmt_3385_sources/type_cast_3391/SplitProtocol/Update/ca
      -- 
    ca_18836_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3391_inst_ack_1, ack => cp_elements(2142)); -- 
    -- CP-element group 2143 join  transition  output  bypass 
    -- predecessors 2140 2142 
    -- successors 2144 
    -- members (6) 
      -- 	branch_block_stmt_2042/xx_xloopexitx_xix_xix_xix_xloopexit_xx_xloopexitx_xix_xix_xi_PhiReq/phi_stmt_3385/phi_stmt_3385_sources/type_cast_3391/SplitProtocol/$exit
      -- 	branch_block_stmt_2042/xx_xloopexitx_xix_xix_xix_xloopexit_xx_xloopexitx_xix_xix_xi_PhiReq/phi_stmt_3385/phi_stmt_3385_sources/type_cast_3391/$exit
      -- 	branch_block_stmt_2042/xx_xloopexitx_xix_xix_xix_xloopexit_xx_xloopexitx_xix_xix_xi_PhiReq/phi_stmt_3385/phi_stmt_3385_sources/$exit
      -- 	branch_block_stmt_2042/xx_xloopexitx_xix_xix_xix_xloopexit_xx_xloopexitx_xix_xix_xi_PhiReq/phi_stmt_3385/$exit
      -- 	branch_block_stmt_2042/xx_xloopexitx_xix_xix_xix_xloopexit_xx_xloopexitx_xix_xix_xi_PhiReq/$exit
      -- 	branch_block_stmt_2042/xx_xloopexitx_xix_xix_xix_xloopexit_xx_xloopexitx_xix_xix_xi_PhiReq/phi_stmt_3385/phi_stmt_3385_req
      -- 
    cp_element_group_2143: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_2143"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(2140) & cp_elements(2142);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(2143), clk => clk, reset => reset); --
    end block;
    phi_stmt_3385_req_18837_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2143), ack => phi_stmt_3385_req_1); -- 
    -- CP-element group 2144 merge  place  bypass 
    -- predecessors 2138 2143 
    -- successors 2145 
    -- members (1) 
      -- 	branch_block_stmt_2042/merge_stmt_3384_PhiReqMerge
      -- 
    cp_elements(2144) <= OrReduce(cp_elements(2138) & cp_elements(2143));
    -- CP-element group 2145 transition  bypass 
    -- predecessors 2144 
    -- successors 2146 
    -- members (1) 
      -- 	branch_block_stmt_2042/merge_stmt_3384_PhiAck/$entry
      -- 
    cp_elements(2145) <= cp_elements(2144);
    -- CP-element group 2146 fork  transition  place  input  bypass 
    -- predecessors 2145 
    -- successors 2158 2164 
    -- members (7) 
      -- 	branch_block_stmt_2042/xx_xloopexitx_xix_xix_xi_udiv32x_xexitx_xpreheaderx_xix_xi
      -- 	branch_block_stmt_2042/merge_stmt_3384__exit__
      -- 	branch_block_stmt_2042/xx_xloopexitx_xix_xix_xi_udiv32x_xexitx_xpreheaderx_xix_xi_PhiReq/phi_stmt_3395/phi_stmt_3395_sources/$entry
      -- 	branch_block_stmt_2042/xx_xloopexitx_xix_xix_xi_udiv32x_xexitx_xpreheaderx_xix_xi_PhiReq/phi_stmt_3395/$entry
      -- 	branch_block_stmt_2042/xx_xloopexitx_xix_xix_xi_udiv32x_xexitx_xpreheaderx_xix_xi_PhiReq/$entry
      -- 	branch_block_stmt_2042/merge_stmt_3384_PhiAck/phi_stmt_3385_ack
      -- 	branch_block_stmt_2042/merge_stmt_3384_PhiAck/$exit
      -- 
    phi_stmt_3385_ack_18842_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_3385_ack_0, ack => cp_elements(2146)); -- 
    -- CP-element group 2147 fork  transition  bypass 
    -- predecessors 824 
    -- successors 2148 2149 
    -- members (2) 
      -- 	branch_block_stmt_2042/bb_41_udiv32x_xexitx_xpreheaderx_xix_xi_PhiReq/phi_stmt_3395/phi_stmt_3395_sources/type_cast_3398/SplitProtocol/$entry
      -- 	branch_block_stmt_2042/bb_41_udiv32x_xexitx_xpreheaderx_xix_xi_PhiReq/phi_stmt_3395/phi_stmt_3395_sources/type_cast_3398/$entry
      -- 
    cp_elements(2147) <= cp_elements(824);
    -- CP-element group 2148 transition  bypass 
    -- predecessors 2147 
    -- successors 2150 
    -- members (4) 
      -- 	branch_block_stmt_2042/bb_41_udiv32x_xexitx_xpreheaderx_xix_xi_PhiReq/phi_stmt_3395/phi_stmt_3395_sources/type_cast_3398/SplitProtocol/Sample/ra
      -- 	branch_block_stmt_2042/bb_41_udiv32x_xexitx_xpreheaderx_xix_xi_PhiReq/phi_stmt_3395/phi_stmt_3395_sources/type_cast_3398/SplitProtocol/Sample/rr
      -- 	branch_block_stmt_2042/bb_41_udiv32x_xexitx_xpreheaderx_xix_xi_PhiReq/phi_stmt_3395/phi_stmt_3395_sources/type_cast_3398/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_2042/bb_41_udiv32x_xexitx_xpreheaderx_xix_xi_PhiReq/phi_stmt_3395/phi_stmt_3395_sources/type_cast_3398/SplitProtocol/Sample/$entry
      -- 
    cp_elements(2148) <= cp_elements(2147);
    -- CP-element group 2149 transition  bypass 
    -- predecessors 2147 
    -- successors 2150 
    -- members (4) 
      -- 	branch_block_stmt_2042/bb_41_udiv32x_xexitx_xpreheaderx_xix_xi_PhiReq/phi_stmt_3395/phi_stmt_3395_sources/type_cast_3398/SplitProtocol/Update/ca
      -- 	branch_block_stmt_2042/bb_41_udiv32x_xexitx_xpreheaderx_xix_xi_PhiReq/phi_stmt_3395/phi_stmt_3395_sources/type_cast_3398/SplitProtocol/Update/cr
      -- 	branch_block_stmt_2042/bb_41_udiv32x_xexitx_xpreheaderx_xix_xi_PhiReq/phi_stmt_3395/phi_stmt_3395_sources/type_cast_3398/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_2042/bb_41_udiv32x_xexitx_xpreheaderx_xix_xi_PhiReq/phi_stmt_3395/phi_stmt_3395_sources/type_cast_3398/SplitProtocol/Update/$entry
      -- 
    cp_elements(2149) <= cp_elements(2147);
    -- CP-element group 2150 join  transition  bypass 
    -- predecessors 2148 2149 
    -- successors 2157 
    -- members (2) 
      -- 	branch_block_stmt_2042/bb_41_udiv32x_xexitx_xpreheaderx_xix_xi_PhiReq/phi_stmt_3395/phi_stmt_3395_sources/type_cast_3398/SplitProtocol/$exit
      -- 	branch_block_stmt_2042/bb_41_udiv32x_xexitx_xpreheaderx_xix_xi_PhiReq/phi_stmt_3395/phi_stmt_3395_sources/type_cast_3398/$exit
      -- 
    cp_element_group_2150: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_2150"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(2148) & cp_elements(2149);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(2150), clk => clk, reset => reset); --
    end block;
    -- CP-element group 2151 fork  transition  bypass 
    -- predecessors 824 
    -- successors 2152 2154 
    -- members (2) 
      -- 	branch_block_stmt_2042/bb_41_udiv32x_xexitx_xpreheaderx_xix_xi_PhiReq/phi_stmt_3395/phi_stmt_3395_sources/type_cast_3400/SplitProtocol/$entry
      -- 	branch_block_stmt_2042/bb_41_udiv32x_xexitx_xpreheaderx_xix_xi_PhiReq/phi_stmt_3395/phi_stmt_3395_sources/type_cast_3400/$entry
      -- 
    cp_elements(2151) <= cp_elements(824);
    -- CP-element group 2152 transition  output  bypass 
    -- predecessors 2151 
    -- successors 2153 
    -- members (2) 
      -- 	branch_block_stmt_2042/bb_41_udiv32x_xexitx_xpreheaderx_xix_xi_PhiReq/phi_stmt_3395/phi_stmt_3395_sources/type_cast_3400/SplitProtocol/Sample/rr
      -- 	branch_block_stmt_2042/bb_41_udiv32x_xexitx_xpreheaderx_xix_xi_PhiReq/phi_stmt_3395/phi_stmt_3395_sources/type_cast_3400/SplitProtocol/Sample/$entry
      -- 
    cp_elements(2152) <= cp_elements(2151);
    rr_18877_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2152), ack => type_cast_3400_inst_req_0); -- 
    -- CP-element group 2153 transition  input  bypass 
    -- predecessors 2152 
    -- successors 2156 
    -- members (2) 
      -- 	branch_block_stmt_2042/bb_41_udiv32x_xexitx_xpreheaderx_xix_xi_PhiReq/phi_stmt_3395/phi_stmt_3395_sources/type_cast_3400/SplitProtocol/Sample/ra
      -- 	branch_block_stmt_2042/bb_41_udiv32x_xexitx_xpreheaderx_xix_xi_PhiReq/phi_stmt_3395/phi_stmt_3395_sources/type_cast_3400/SplitProtocol/Sample/$exit
      -- 
    ra_18878_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3400_inst_ack_0, ack => cp_elements(2153)); -- 
    -- CP-element group 2154 transition  output  bypass 
    -- predecessors 2151 
    -- successors 2155 
    -- members (2) 
      -- 	branch_block_stmt_2042/bb_41_udiv32x_xexitx_xpreheaderx_xix_xi_PhiReq/phi_stmt_3395/phi_stmt_3395_sources/type_cast_3400/SplitProtocol/Update/cr
      -- 	branch_block_stmt_2042/bb_41_udiv32x_xexitx_xpreheaderx_xix_xi_PhiReq/phi_stmt_3395/phi_stmt_3395_sources/type_cast_3400/SplitProtocol/Update/$entry
      -- 
    cp_elements(2154) <= cp_elements(2151);
    cr_18882_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2154), ack => type_cast_3400_inst_req_1); -- 
    -- CP-element group 2155 transition  input  bypass 
    -- predecessors 2154 
    -- successors 2156 
    -- members (2) 
      -- 	branch_block_stmt_2042/bb_41_udiv32x_xexitx_xpreheaderx_xix_xi_PhiReq/phi_stmt_3395/phi_stmt_3395_sources/type_cast_3400/SplitProtocol/Update/ca
      -- 	branch_block_stmt_2042/bb_41_udiv32x_xexitx_xpreheaderx_xix_xi_PhiReq/phi_stmt_3395/phi_stmt_3395_sources/type_cast_3400/SplitProtocol/Update/$exit
      -- 
    ca_18883_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3400_inst_ack_1, ack => cp_elements(2155)); -- 
    -- CP-element group 2156 join  transition  bypass 
    -- predecessors 2153 2155 
    -- successors 2157 
    -- members (2) 
      -- 	branch_block_stmt_2042/bb_41_udiv32x_xexitx_xpreheaderx_xix_xi_PhiReq/phi_stmt_3395/phi_stmt_3395_sources/type_cast_3400/SplitProtocol/$exit
      -- 	branch_block_stmt_2042/bb_41_udiv32x_xexitx_xpreheaderx_xix_xi_PhiReq/phi_stmt_3395/phi_stmt_3395_sources/type_cast_3400/$exit
      -- 
    cp_element_group_2156: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_2156"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(2153) & cp_elements(2155);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(2156), clk => clk, reset => reset); --
    end block;
    -- CP-element group 2157 join  transition  output  bypass 
    -- predecessors 2150 2156 
    -- successors 2169 
    -- members (4) 
      -- 	branch_block_stmt_2042/bb_41_udiv32x_xexitx_xpreheaderx_xix_xi_PhiReq/phi_stmt_3395/phi_stmt_3395_req
      -- 	branch_block_stmt_2042/bb_41_udiv32x_xexitx_xpreheaderx_xix_xi_PhiReq/phi_stmt_3395/phi_stmt_3395_sources/$exit
      -- 	branch_block_stmt_2042/bb_41_udiv32x_xexitx_xpreheaderx_xix_xi_PhiReq/phi_stmt_3395/$exit
      -- 	branch_block_stmt_2042/bb_41_udiv32x_xexitx_xpreheaderx_xix_xi_PhiReq/$exit
      -- 
    cp_element_group_2157: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_2157"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(2150) & cp_elements(2156);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(2157), clk => clk, reset => reset); --
    end block;
    phi_stmt_3395_req_18884_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2157), ack => phi_stmt_3395_req_1); -- 
    -- CP-element group 2158 fork  transition  bypass 
    -- predecessors 2146 
    -- successors 2159 2161 
    -- members (2) 
      -- 	branch_block_stmt_2042/xx_xloopexitx_xix_xix_xi_udiv32x_xexitx_xpreheaderx_xix_xi_PhiReq/phi_stmt_3395/phi_stmt_3395_sources/type_cast_3398/SplitProtocol/$entry
      -- 	branch_block_stmt_2042/xx_xloopexitx_xix_xix_xi_udiv32x_xexitx_xpreheaderx_xix_xi_PhiReq/phi_stmt_3395/phi_stmt_3395_sources/type_cast_3398/$entry
      -- 
    cp_elements(2158) <= cp_elements(2146);
    -- CP-element group 2159 transition  output  bypass 
    -- predecessors 2158 
    -- successors 2160 
    -- members (2) 
      -- 	branch_block_stmt_2042/xx_xloopexitx_xix_xix_xi_udiv32x_xexitx_xpreheaderx_xix_xi_PhiReq/phi_stmt_3395/phi_stmt_3395_sources/type_cast_3398/SplitProtocol/Sample/rr
      -- 	branch_block_stmt_2042/xx_xloopexitx_xix_xix_xi_udiv32x_xexitx_xpreheaderx_xix_xi_PhiReq/phi_stmt_3395/phi_stmt_3395_sources/type_cast_3398/SplitProtocol/Sample/$entry
      -- 
    cp_elements(2159) <= cp_elements(2158);
    rr_18903_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2159), ack => type_cast_3398_inst_req_0); -- 
    -- CP-element group 2160 transition  input  bypass 
    -- predecessors 2159 
    -- successors 2163 
    -- members (2) 
      -- 	branch_block_stmt_2042/xx_xloopexitx_xix_xix_xi_udiv32x_xexitx_xpreheaderx_xix_xi_PhiReq/phi_stmt_3395/phi_stmt_3395_sources/type_cast_3398/SplitProtocol/Sample/ra
      -- 	branch_block_stmt_2042/xx_xloopexitx_xix_xix_xi_udiv32x_xexitx_xpreheaderx_xix_xi_PhiReq/phi_stmt_3395/phi_stmt_3395_sources/type_cast_3398/SplitProtocol/Sample/$exit
      -- 
    ra_18904_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3398_inst_ack_0, ack => cp_elements(2160)); -- 
    -- CP-element group 2161 transition  output  bypass 
    -- predecessors 2158 
    -- successors 2162 
    -- members (2) 
      -- 	branch_block_stmt_2042/xx_xloopexitx_xix_xix_xi_udiv32x_xexitx_xpreheaderx_xix_xi_PhiReq/phi_stmt_3395/phi_stmt_3395_sources/type_cast_3398/SplitProtocol/Update/cr
      -- 	branch_block_stmt_2042/xx_xloopexitx_xix_xix_xi_udiv32x_xexitx_xpreheaderx_xix_xi_PhiReq/phi_stmt_3395/phi_stmt_3395_sources/type_cast_3398/SplitProtocol/Update/$entry
      -- 
    cp_elements(2161) <= cp_elements(2158);
    cr_18908_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2161), ack => type_cast_3398_inst_req_1); -- 
    -- CP-element group 2162 transition  input  bypass 
    -- predecessors 2161 
    -- successors 2163 
    -- members (2) 
      -- 	branch_block_stmt_2042/xx_xloopexitx_xix_xix_xi_udiv32x_xexitx_xpreheaderx_xix_xi_PhiReq/phi_stmt_3395/phi_stmt_3395_sources/type_cast_3398/SplitProtocol/Update/ca
      -- 	branch_block_stmt_2042/xx_xloopexitx_xix_xix_xi_udiv32x_xexitx_xpreheaderx_xix_xi_PhiReq/phi_stmt_3395/phi_stmt_3395_sources/type_cast_3398/SplitProtocol/Update/$exit
      -- 
    ca_18909_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3398_inst_ack_1, ack => cp_elements(2162)); -- 
    -- CP-element group 2163 join  transition  bypass 
    -- predecessors 2160 2162 
    -- successors 2168 
    -- members (2) 
      -- 	branch_block_stmt_2042/xx_xloopexitx_xix_xix_xi_udiv32x_xexitx_xpreheaderx_xix_xi_PhiReq/phi_stmt_3395/phi_stmt_3395_sources/type_cast_3398/SplitProtocol/$exit
      -- 	branch_block_stmt_2042/xx_xloopexitx_xix_xix_xi_udiv32x_xexitx_xpreheaderx_xix_xi_PhiReq/phi_stmt_3395/phi_stmt_3395_sources/type_cast_3398/$exit
      -- 
    cp_element_group_2163: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_2163"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(2160) & cp_elements(2162);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(2163), clk => clk, reset => reset); --
    end block;
    -- CP-element group 2164 fork  transition  bypass 
    -- predecessors 2146 
    -- successors 2165 2166 
    -- members (2) 
      -- 	branch_block_stmt_2042/xx_xloopexitx_xix_xix_xi_udiv32x_xexitx_xpreheaderx_xix_xi_PhiReq/phi_stmt_3395/phi_stmt_3395_sources/type_cast_3400/SplitProtocol/$entry
      -- 	branch_block_stmt_2042/xx_xloopexitx_xix_xix_xi_udiv32x_xexitx_xpreheaderx_xix_xi_PhiReq/phi_stmt_3395/phi_stmt_3395_sources/type_cast_3400/$entry
      -- 
    cp_elements(2164) <= cp_elements(2146);
    -- CP-element group 2165 transition  bypass 
    -- predecessors 2164 
    -- successors 2167 
    -- members (4) 
      -- 	branch_block_stmt_2042/xx_xloopexitx_xix_xix_xi_udiv32x_xexitx_xpreheaderx_xix_xi_PhiReq/phi_stmt_3395/phi_stmt_3395_sources/type_cast_3400/SplitProtocol/Sample/ra
      -- 	branch_block_stmt_2042/xx_xloopexitx_xix_xix_xi_udiv32x_xexitx_xpreheaderx_xix_xi_PhiReq/phi_stmt_3395/phi_stmt_3395_sources/type_cast_3400/SplitProtocol/Sample/rr
      -- 	branch_block_stmt_2042/xx_xloopexitx_xix_xix_xi_udiv32x_xexitx_xpreheaderx_xix_xi_PhiReq/phi_stmt_3395/phi_stmt_3395_sources/type_cast_3400/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_2042/xx_xloopexitx_xix_xix_xi_udiv32x_xexitx_xpreheaderx_xix_xi_PhiReq/phi_stmt_3395/phi_stmt_3395_sources/type_cast_3400/SplitProtocol/Sample/$entry
      -- 
    cp_elements(2165) <= cp_elements(2164);
    -- CP-element group 2166 transition  bypass 
    -- predecessors 2164 
    -- successors 2167 
    -- members (4) 
      -- 	branch_block_stmt_2042/xx_xloopexitx_xix_xix_xi_udiv32x_xexitx_xpreheaderx_xix_xi_PhiReq/phi_stmt_3395/phi_stmt_3395_sources/type_cast_3400/SplitProtocol/Update/ca
      -- 	branch_block_stmt_2042/xx_xloopexitx_xix_xix_xi_udiv32x_xexitx_xpreheaderx_xix_xi_PhiReq/phi_stmt_3395/phi_stmt_3395_sources/type_cast_3400/SplitProtocol/Update/cr
      -- 	branch_block_stmt_2042/xx_xloopexitx_xix_xix_xi_udiv32x_xexitx_xpreheaderx_xix_xi_PhiReq/phi_stmt_3395/phi_stmt_3395_sources/type_cast_3400/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_2042/xx_xloopexitx_xix_xix_xi_udiv32x_xexitx_xpreheaderx_xix_xi_PhiReq/phi_stmt_3395/phi_stmt_3395_sources/type_cast_3400/SplitProtocol/Update/$entry
      -- 
    cp_elements(2166) <= cp_elements(2164);
    -- CP-element group 2167 join  transition  bypass 
    -- predecessors 2165 2166 
    -- successors 2168 
    -- members (2) 
      -- 	branch_block_stmt_2042/xx_xloopexitx_xix_xix_xi_udiv32x_xexitx_xpreheaderx_xix_xi_PhiReq/phi_stmt_3395/phi_stmt_3395_sources/type_cast_3400/SplitProtocol/$exit
      -- 	branch_block_stmt_2042/xx_xloopexitx_xix_xix_xi_udiv32x_xexitx_xpreheaderx_xix_xi_PhiReq/phi_stmt_3395/phi_stmt_3395_sources/type_cast_3400/$exit
      -- 
    cp_element_group_2167: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_2167"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(2165) & cp_elements(2166);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(2167), clk => clk, reset => reset); --
    end block;
    -- CP-element group 2168 join  transition  output  bypass 
    -- predecessors 2163 2167 
    -- successors 2169 
    -- members (4) 
      -- 	branch_block_stmt_2042/xx_xloopexitx_xix_xix_xi_udiv32x_xexitx_xpreheaderx_xix_xi_PhiReq/phi_stmt_3395/phi_stmt_3395_req
      -- 	branch_block_stmt_2042/xx_xloopexitx_xix_xix_xi_udiv32x_xexitx_xpreheaderx_xix_xi_PhiReq/phi_stmt_3395/phi_stmt_3395_sources/$exit
      -- 	branch_block_stmt_2042/xx_xloopexitx_xix_xix_xi_udiv32x_xexitx_xpreheaderx_xix_xi_PhiReq/phi_stmt_3395/$exit
      -- 	branch_block_stmt_2042/xx_xloopexitx_xix_xix_xi_udiv32x_xexitx_xpreheaderx_xix_xi_PhiReq/$exit
      -- 
    cp_element_group_2168: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_2168"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(2163) & cp_elements(2167);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(2168), clk => clk, reset => reset); --
    end block;
    phi_stmt_3395_req_18926_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2168), ack => phi_stmt_3395_req_0); -- 
    -- CP-element group 2169 merge  place  bypass 
    -- predecessors 2157 2168 
    -- successors 2170 
    -- members (1) 
      -- 	branch_block_stmt_2042/merge_stmt_3394_PhiReqMerge
      -- 
    cp_elements(2169) <= OrReduce(cp_elements(2157) & cp_elements(2168));
    -- CP-element group 2170 transition  bypass 
    -- predecessors 2169 
    -- successors 2171 
    -- members (1) 
      -- 	branch_block_stmt_2042/merge_stmt_3394_PhiAck/$entry
      -- 
    cp_elements(2170) <= cp_elements(2169);
    -- CP-element group 2171 transition  place  input  bypass 
    -- predecessors 2170 
    -- successors 892 
    -- members (4) 
      -- 	branch_block_stmt_2042/assign_stmt_3407_to_assign_stmt_3426__entry__
      -- 	branch_block_stmt_2042/merge_stmt_3394__exit__
      -- 	branch_block_stmt_2042/merge_stmt_3394_PhiAck/phi_stmt_3395_ack
      -- 	branch_block_stmt_2042/merge_stmt_3394_PhiAck/$exit
      -- 
    phi_stmt_3395_ack_18931_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_3395_ack_0, ack => cp_elements(2171)); -- 
    -- CP-element group 2172 fork  transition  bypass 
    -- predecessors 948 
    -- successors 2173 2185 
    -- members (1) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi_udiv32x_xexitx_xix_xi_PhiReq/$entry
      -- 
    cp_elements(2172) <= cp_elements(948);
    -- CP-element group 2173 fork  transition  bypass 
    -- predecessors 2172 
    -- successors 2174 2180 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi_udiv32x_xexitx_xix_xi_PhiReq/phi_stmt_3443/phi_stmt_3443_sources/$entry
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi_udiv32x_xexitx_xix_xi_PhiReq/phi_stmt_3443/$entry
      -- 
    cp_elements(2173) <= cp_elements(2172);
    -- CP-element group 2174 fork  transition  bypass 
    -- predecessors 2173 
    -- successors 2175 2177 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi_udiv32x_xexitx_xix_xi_PhiReq/phi_stmt_3443/phi_stmt_3443_sources/type_cast_3446/$entry
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi_udiv32x_xexitx_xix_xi_PhiReq/phi_stmt_3443/phi_stmt_3443_sources/type_cast_3446/SplitProtocol/$entry
      -- 
    cp_elements(2174) <= cp_elements(2173);
    -- CP-element group 2175 transition  output  bypass 
    -- predecessors 2174 
    -- successors 2176 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi_udiv32x_xexitx_xix_xi_PhiReq/phi_stmt_3443/phi_stmt_3443_sources/type_cast_3446/SplitProtocol/Sample/rr
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi_udiv32x_xexitx_xix_xi_PhiReq/phi_stmt_3443/phi_stmt_3443_sources/type_cast_3446/SplitProtocol/Sample/$entry
      -- 
    cp_elements(2175) <= cp_elements(2174);
    rr_18962_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2175), ack => type_cast_3446_inst_req_0); -- 
    -- CP-element group 2176 transition  input  bypass 
    -- predecessors 2175 
    -- successors 2179 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi_udiv32x_xexitx_xix_xi_PhiReq/phi_stmt_3443/phi_stmt_3443_sources/type_cast_3446/SplitProtocol/Sample/ra
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi_udiv32x_xexitx_xix_xi_PhiReq/phi_stmt_3443/phi_stmt_3443_sources/type_cast_3446/SplitProtocol/Sample/$exit
      -- 
    ra_18963_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3446_inst_ack_0, ack => cp_elements(2176)); -- 
    -- CP-element group 2177 transition  output  bypass 
    -- predecessors 2174 
    -- successors 2178 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi_udiv32x_xexitx_xix_xi_PhiReq/phi_stmt_3443/phi_stmt_3443_sources/type_cast_3446/SplitProtocol/Update/cr
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi_udiv32x_xexitx_xix_xi_PhiReq/phi_stmt_3443/phi_stmt_3443_sources/type_cast_3446/SplitProtocol/Update/$entry
      -- 
    cp_elements(2177) <= cp_elements(2174);
    cr_18967_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2177), ack => type_cast_3446_inst_req_1); -- 
    -- CP-element group 2178 transition  input  bypass 
    -- predecessors 2177 
    -- successors 2179 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi_udiv32x_xexitx_xix_xi_PhiReq/phi_stmt_3443/phi_stmt_3443_sources/type_cast_3446/SplitProtocol/Update/ca
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi_udiv32x_xexitx_xix_xi_PhiReq/phi_stmt_3443/phi_stmt_3443_sources/type_cast_3446/SplitProtocol/Update/$exit
      -- 
    ca_18968_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3446_inst_ack_1, ack => cp_elements(2178)); -- 
    -- CP-element group 2179 join  transition  bypass 
    -- predecessors 2176 2178 
    -- successors 2184 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi_udiv32x_xexitx_xix_xi_PhiReq/phi_stmt_3443/phi_stmt_3443_sources/type_cast_3446/SplitProtocol/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi_udiv32x_xexitx_xix_xi_PhiReq/phi_stmt_3443/phi_stmt_3443_sources/type_cast_3446/$exit
      -- 
    cp_element_group_2179: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_2179"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(2176) & cp_elements(2178);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(2179), clk => clk, reset => reset); --
    end block;
    -- CP-element group 2180 fork  transition  bypass 
    -- predecessors 2173 
    -- successors 2181 2182 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi_udiv32x_xexitx_xix_xi_PhiReq/phi_stmt_3443/phi_stmt_3443_sources/type_cast_3448/$entry
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi_udiv32x_xexitx_xix_xi_PhiReq/phi_stmt_3443/phi_stmt_3443_sources/type_cast_3448/SplitProtocol/$entry
      -- 
    cp_elements(2180) <= cp_elements(2173);
    -- CP-element group 2181 transition  bypass 
    -- predecessors 2180 
    -- successors 2183 
    -- members (4) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi_udiv32x_xexitx_xix_xi_PhiReq/phi_stmt_3443/phi_stmt_3443_sources/type_cast_3448/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi_udiv32x_xexitx_xix_xi_PhiReq/phi_stmt_3443/phi_stmt_3443_sources/type_cast_3448/SplitProtocol/Sample/rr
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi_udiv32x_xexitx_xix_xi_PhiReq/phi_stmt_3443/phi_stmt_3443_sources/type_cast_3448/SplitProtocol/Sample/ra
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi_udiv32x_xexitx_xix_xi_PhiReq/phi_stmt_3443/phi_stmt_3443_sources/type_cast_3448/SplitProtocol/Sample/$entry
      -- 
    cp_elements(2181) <= cp_elements(2180);
    -- CP-element group 2182 transition  bypass 
    -- predecessors 2180 
    -- successors 2183 
    -- members (4) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi_udiv32x_xexitx_xix_xi_PhiReq/phi_stmt_3443/phi_stmt_3443_sources/type_cast_3448/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi_udiv32x_xexitx_xix_xi_PhiReq/phi_stmt_3443/phi_stmt_3443_sources/type_cast_3448/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi_udiv32x_xexitx_xix_xi_PhiReq/phi_stmt_3443/phi_stmt_3443_sources/type_cast_3448/SplitProtocol/Update/cr
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi_udiv32x_xexitx_xix_xi_PhiReq/phi_stmt_3443/phi_stmt_3443_sources/type_cast_3448/SplitProtocol/Update/ca
      -- 
    cp_elements(2182) <= cp_elements(2180);
    -- CP-element group 2183 join  transition  bypass 
    -- predecessors 2181 2182 
    -- successors 2184 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi_udiv32x_xexitx_xix_xi_PhiReq/phi_stmt_3443/phi_stmt_3443_sources/type_cast_3448/SplitProtocol/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi_udiv32x_xexitx_xix_xi_PhiReq/phi_stmt_3443/phi_stmt_3443_sources/type_cast_3448/$exit
      -- 
    cp_element_group_2183: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_2183"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(2181) & cp_elements(2182);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(2183), clk => clk, reset => reset); --
    end block;
    -- CP-element group 2184 join  transition  output  bypass 
    -- predecessors 2179 2183 
    -- successors 2191 
    -- members (3) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi_udiv32x_xexitx_xix_xi_PhiReq/phi_stmt_3443/phi_stmt_3443_req
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi_udiv32x_xexitx_xix_xi_PhiReq/phi_stmt_3443/phi_stmt_3443_sources/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi_udiv32x_xexitx_xix_xi_PhiReq/phi_stmt_3443/$exit
      -- 
    cp_element_group_2184: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_2184"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(2179) & cp_elements(2183);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(2184), clk => clk, reset => reset); --
    end block;
    phi_stmt_3443_req_18985_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2184), ack => phi_stmt_3443_req_0); -- 
    -- CP-element group 2185 fork  transition  bypass 
    -- predecessors 2172 
    -- successors 2186 2188 
    -- members (4) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi_udiv32x_xexitx_xix_xi_PhiReq/phi_stmt_3436/phi_stmt_3436_sources/$entry
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi_udiv32x_xexitx_xix_xi_PhiReq/phi_stmt_3436/$entry
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi_udiv32x_xexitx_xix_xi_PhiReq/phi_stmt_3436/phi_stmt_3436_sources/type_cast_3439/SplitProtocol/$entry
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi_udiv32x_xexitx_xix_xi_PhiReq/phi_stmt_3436/phi_stmt_3436_sources/type_cast_3439/$entry
      -- 
    cp_elements(2185) <= cp_elements(2172);
    -- CP-element group 2186 transition  output  bypass 
    -- predecessors 2185 
    -- successors 2187 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi_udiv32x_xexitx_xix_xi_PhiReq/phi_stmt_3436/phi_stmt_3436_sources/type_cast_3439/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi_udiv32x_xexitx_xix_xi_PhiReq/phi_stmt_3436/phi_stmt_3436_sources/type_cast_3439/SplitProtocol/Sample/rr
      -- 
    cp_elements(2186) <= cp_elements(2185);
    rr_19001_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2186), ack => type_cast_3439_inst_req_0); -- 
    -- CP-element group 2187 transition  input  bypass 
    -- predecessors 2186 
    -- successors 2190 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi_udiv32x_xexitx_xix_xi_PhiReq/phi_stmt_3436/phi_stmt_3436_sources/type_cast_3439/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi_udiv32x_xexitx_xix_xi_PhiReq/phi_stmt_3436/phi_stmt_3436_sources/type_cast_3439/SplitProtocol/Sample/ra
      -- 
    ra_19002_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3439_inst_ack_0, ack => cp_elements(2187)); -- 
    -- CP-element group 2188 transition  output  bypass 
    -- predecessors 2185 
    -- successors 2189 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi_udiv32x_xexitx_xix_xi_PhiReq/phi_stmt_3436/phi_stmt_3436_sources/type_cast_3439/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi_udiv32x_xexitx_xix_xi_PhiReq/phi_stmt_3436/phi_stmt_3436_sources/type_cast_3439/SplitProtocol/Update/cr
      -- 
    cp_elements(2188) <= cp_elements(2185);
    cr_19006_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2188), ack => type_cast_3439_inst_req_1); -- 
    -- CP-element group 2189 transition  input  bypass 
    -- predecessors 2188 
    -- successors 2190 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi_udiv32x_xexitx_xix_xi_PhiReq/phi_stmt_3436/phi_stmt_3436_sources/type_cast_3439/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi_udiv32x_xexitx_xix_xi_PhiReq/phi_stmt_3436/phi_stmt_3436_sources/type_cast_3439/SplitProtocol/Update/ca
      -- 
    ca_19007_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3439_inst_ack_1, ack => cp_elements(2189)); -- 
    -- CP-element group 2190 join  transition  output  bypass 
    -- predecessors 2187 2189 
    -- successors 2191 
    -- members (5) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi_udiv32x_xexitx_xix_xi_PhiReq/phi_stmt_3436/phi_stmt_3436_sources/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi_udiv32x_xexitx_xix_xi_PhiReq/phi_stmt_3436/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi_udiv32x_xexitx_xix_xi_PhiReq/phi_stmt_3436/phi_stmt_3436_sources/type_cast_3439/SplitProtocol/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi_udiv32x_xexitx_xix_xi_PhiReq/phi_stmt_3436/phi_stmt_3436_sources/type_cast_3439/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi_udiv32x_xexitx_xix_xi_PhiReq/phi_stmt_3436/phi_stmt_3436_req
      -- 
    cp_element_group_2190: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_2190"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(2187) & cp_elements(2189);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(2190), clk => clk, reset => reset); --
    end block;
    phi_stmt_3436_req_19008_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2190), ack => phi_stmt_3436_req_0); -- 
    -- CP-element group 2191 join  transition  bypass 
    -- predecessors 2184 2190 
    -- successors 2210 
    -- members (1) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi_udiv32x_xexitx_xix_xi_PhiReq/$exit
      -- 
    cp_element_group_2191: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_2191"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(2184) & cp_elements(2190);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(2191), clk => clk, reset => reset); --
    end block;
    -- CP-element group 2192 fork  transition  bypass 
    -- predecessors 55 
    -- successors 2193 2205 
    -- members (1) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xix_xpreheader_udiv32x_xexitx_xix_xi_PhiReq/$entry
      -- 
    cp_elements(2192) <= cp_elements(55);
    -- CP-element group 2193 fork  transition  bypass 
    -- predecessors 2192 
    -- successors 2194 2198 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xix_xpreheader_udiv32x_xexitx_xix_xi_PhiReq/phi_stmt_3443/$entry
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xix_xpreheader_udiv32x_xexitx_xix_xi_PhiReq/phi_stmt_3443/phi_stmt_3443_sources/$entry
      -- 
    cp_elements(2193) <= cp_elements(2192);
    -- CP-element group 2194 fork  transition  bypass 
    -- predecessors 2193 
    -- successors 2195 2196 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xix_xpreheader_udiv32x_xexitx_xix_xi_PhiReq/phi_stmt_3443/phi_stmt_3443_sources/type_cast_3446/$entry
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xix_xpreheader_udiv32x_xexitx_xix_xi_PhiReq/phi_stmt_3443/phi_stmt_3443_sources/type_cast_3446/SplitProtocol/$entry
      -- 
    cp_elements(2194) <= cp_elements(2193);
    -- CP-element group 2195 transition  bypass 
    -- predecessors 2194 
    -- successors 2197 
    -- members (4) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xix_xpreheader_udiv32x_xexitx_xix_xi_PhiReq/phi_stmt_3443/phi_stmt_3443_sources/type_cast_3446/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xix_xpreheader_udiv32x_xexitx_xix_xi_PhiReq/phi_stmt_3443/phi_stmt_3443_sources/type_cast_3446/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xix_xpreheader_udiv32x_xexitx_xix_xi_PhiReq/phi_stmt_3443/phi_stmt_3443_sources/type_cast_3446/SplitProtocol/Sample/rr
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xix_xpreheader_udiv32x_xexitx_xix_xi_PhiReq/phi_stmt_3443/phi_stmt_3443_sources/type_cast_3446/SplitProtocol/Sample/ra
      -- 
    cp_elements(2195) <= cp_elements(2194);
    -- CP-element group 2196 transition  bypass 
    -- predecessors 2194 
    -- successors 2197 
    -- members (4) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xix_xpreheader_udiv32x_xexitx_xix_xi_PhiReq/phi_stmt_3443/phi_stmt_3443_sources/type_cast_3446/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xix_xpreheader_udiv32x_xexitx_xix_xi_PhiReq/phi_stmt_3443/phi_stmt_3443_sources/type_cast_3446/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xix_xpreheader_udiv32x_xexitx_xix_xi_PhiReq/phi_stmt_3443/phi_stmt_3443_sources/type_cast_3446/SplitProtocol/Update/cr
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xix_xpreheader_udiv32x_xexitx_xix_xi_PhiReq/phi_stmt_3443/phi_stmt_3443_sources/type_cast_3446/SplitProtocol/Update/ca
      -- 
    cp_elements(2196) <= cp_elements(2194);
    -- CP-element group 2197 join  transition  bypass 
    -- predecessors 2195 2196 
    -- successors 2204 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xix_xpreheader_udiv32x_xexitx_xix_xi_PhiReq/phi_stmt_3443/phi_stmt_3443_sources/type_cast_3446/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xix_xpreheader_udiv32x_xexitx_xix_xi_PhiReq/phi_stmt_3443/phi_stmt_3443_sources/type_cast_3446/SplitProtocol/$exit
      -- 
    cp_element_group_2197: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_2197"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(2195) & cp_elements(2196);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(2197), clk => clk, reset => reset); --
    end block;
    -- CP-element group 2198 fork  transition  bypass 
    -- predecessors 2193 
    -- successors 2199 2201 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xix_xpreheader_udiv32x_xexitx_xix_xi_PhiReq/phi_stmt_3443/phi_stmt_3443_sources/type_cast_3448/$entry
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xix_xpreheader_udiv32x_xexitx_xix_xi_PhiReq/phi_stmt_3443/phi_stmt_3443_sources/type_cast_3448/SplitProtocol/$entry
      -- 
    cp_elements(2198) <= cp_elements(2193);
    -- CP-element group 2199 transition  output  bypass 
    -- predecessors 2198 
    -- successors 2200 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xix_xpreheader_udiv32x_xexitx_xix_xi_PhiReq/phi_stmt_3443/phi_stmt_3443_sources/type_cast_3448/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xix_xpreheader_udiv32x_xexitx_xix_xi_PhiReq/phi_stmt_3443/phi_stmt_3443_sources/type_cast_3448/SplitProtocol/Sample/rr
      -- 
    cp_elements(2199) <= cp_elements(2198);
    rr_19043_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2199), ack => type_cast_3448_inst_req_0); -- 
    -- CP-element group 2200 transition  input  bypass 
    -- predecessors 2199 
    -- successors 2203 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xix_xpreheader_udiv32x_xexitx_xix_xi_PhiReq/phi_stmt_3443/phi_stmt_3443_sources/type_cast_3448/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xix_xpreheader_udiv32x_xexitx_xix_xi_PhiReq/phi_stmt_3443/phi_stmt_3443_sources/type_cast_3448/SplitProtocol/Sample/ra
      -- 
    ra_19044_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3448_inst_ack_0, ack => cp_elements(2200)); -- 
    -- CP-element group 2201 transition  output  bypass 
    -- predecessors 2198 
    -- successors 2202 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xix_xpreheader_udiv32x_xexitx_xix_xi_PhiReq/phi_stmt_3443/phi_stmt_3443_sources/type_cast_3448/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xix_xpreheader_udiv32x_xexitx_xix_xi_PhiReq/phi_stmt_3443/phi_stmt_3443_sources/type_cast_3448/SplitProtocol/Update/cr
      -- 
    cp_elements(2201) <= cp_elements(2198);
    cr_19048_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2201), ack => type_cast_3448_inst_req_1); -- 
    -- CP-element group 2202 transition  input  bypass 
    -- predecessors 2201 
    -- successors 2203 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xix_xpreheader_udiv32x_xexitx_xix_xi_PhiReq/phi_stmt_3443/phi_stmt_3443_sources/type_cast_3448/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xix_xpreheader_udiv32x_xexitx_xix_xi_PhiReq/phi_stmt_3443/phi_stmt_3443_sources/type_cast_3448/SplitProtocol/Update/ca
      -- 
    ca_19049_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3448_inst_ack_1, ack => cp_elements(2202)); -- 
    -- CP-element group 2203 join  transition  bypass 
    -- predecessors 2200 2202 
    -- successors 2204 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xix_xpreheader_udiv32x_xexitx_xix_xi_PhiReq/phi_stmt_3443/phi_stmt_3443_sources/type_cast_3448/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xix_xpreheader_udiv32x_xexitx_xix_xi_PhiReq/phi_stmt_3443/phi_stmt_3443_sources/type_cast_3448/SplitProtocol/$exit
      -- 
    cp_element_group_2203: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_2203"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(2200) & cp_elements(2202);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(2203), clk => clk, reset => reset); --
    end block;
    -- CP-element group 2204 join  transition  output  bypass 
    -- predecessors 2197 2203 
    -- successors 2209 
    -- members (3) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xix_xpreheader_udiv32x_xexitx_xix_xi_PhiReq/phi_stmt_3443/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xix_xpreheader_udiv32x_xexitx_xix_xi_PhiReq/phi_stmt_3443/phi_stmt_3443_sources/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xix_xpreheader_udiv32x_xexitx_xix_xi_PhiReq/phi_stmt_3443/phi_stmt_3443_req
      -- 
    cp_element_group_2204: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_2204"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(2197) & cp_elements(2203);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(2204), clk => clk, reset => reset); --
    end block;
    phi_stmt_3443_req_19050_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2204), ack => phi_stmt_3443_req_1); -- 
    -- CP-element group 2205 fork  transition  bypass 
    -- predecessors 2192 
    -- successors 2206 2207 
    -- members (4) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xix_xpreheader_udiv32x_xexitx_xix_xi_PhiReq/phi_stmt_3436/$entry
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xix_xpreheader_udiv32x_xexitx_xix_xi_PhiReq/phi_stmt_3436/phi_stmt_3436_sources/$entry
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xix_xpreheader_udiv32x_xexitx_xix_xi_PhiReq/phi_stmt_3436/phi_stmt_3436_sources/type_cast_3439/$entry
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xix_xpreheader_udiv32x_xexitx_xix_xi_PhiReq/phi_stmt_3436/phi_stmt_3436_sources/type_cast_3439/SplitProtocol/$entry
      -- 
    cp_elements(2205) <= cp_elements(2192);
    -- CP-element group 2206 transition  bypass 
    -- predecessors 2205 
    -- successors 2208 
    -- members (4) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xix_xpreheader_udiv32x_xexitx_xix_xi_PhiReq/phi_stmt_3436/phi_stmt_3436_sources/type_cast_3439/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xix_xpreheader_udiv32x_xexitx_xix_xi_PhiReq/phi_stmt_3436/phi_stmt_3436_sources/type_cast_3439/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xix_xpreheader_udiv32x_xexitx_xix_xi_PhiReq/phi_stmt_3436/phi_stmt_3436_sources/type_cast_3439/SplitProtocol/Sample/rr
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xix_xpreheader_udiv32x_xexitx_xix_xi_PhiReq/phi_stmt_3436/phi_stmt_3436_sources/type_cast_3439/SplitProtocol/Sample/ra
      -- 
    cp_elements(2206) <= cp_elements(2205);
    -- CP-element group 2207 transition  bypass 
    -- predecessors 2205 
    -- successors 2208 
    -- members (4) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xix_xpreheader_udiv32x_xexitx_xix_xi_PhiReq/phi_stmt_3436/phi_stmt_3436_sources/type_cast_3439/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xix_xpreheader_udiv32x_xexitx_xix_xi_PhiReq/phi_stmt_3436/phi_stmt_3436_sources/type_cast_3439/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xix_xpreheader_udiv32x_xexitx_xix_xi_PhiReq/phi_stmt_3436/phi_stmt_3436_sources/type_cast_3439/SplitProtocol/Update/cr
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xix_xpreheader_udiv32x_xexitx_xix_xi_PhiReq/phi_stmt_3436/phi_stmt_3436_sources/type_cast_3439/SplitProtocol/Update/ca
      -- 
    cp_elements(2207) <= cp_elements(2205);
    -- CP-element group 2208 join  transition  output  bypass 
    -- predecessors 2206 2207 
    -- successors 2209 
    -- members (5) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xix_xpreheader_udiv32x_xexitx_xix_xi_PhiReq/phi_stmt_3436/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xix_xpreheader_udiv32x_xexitx_xix_xi_PhiReq/phi_stmt_3436/phi_stmt_3436_sources/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xix_xpreheader_udiv32x_xexitx_xix_xi_PhiReq/phi_stmt_3436/phi_stmt_3436_sources/type_cast_3439/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xix_xpreheader_udiv32x_xexitx_xix_xi_PhiReq/phi_stmt_3436/phi_stmt_3436_sources/type_cast_3439/SplitProtocol/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xix_xpreheader_udiv32x_xexitx_xix_xi_PhiReq/phi_stmt_3436/phi_stmt_3436_req
      -- 
    cp_element_group_2208: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_2208"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(2206) & cp_elements(2207);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(2208), clk => clk, reset => reset); --
    end block;
    phi_stmt_3436_req_19073_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2208), ack => phi_stmt_3436_req_1); -- 
    -- CP-element group 2209 join  transition  bypass 
    -- predecessors 2204 2208 
    -- successors 2210 
    -- members (1) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xix_xpreheader_udiv32x_xexitx_xix_xi_PhiReq/$exit
      -- 
    cp_element_group_2209: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_2209"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(2204) & cp_elements(2208);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(2209), clk => clk, reset => reset); --
    end block;
    -- CP-element group 2210 merge  place  bypass 
    -- predecessors 2191 2209 
    -- successors 2211 
    -- members (1) 
      -- 	branch_block_stmt_2042/merge_stmt_3435_PhiReqMerge
      -- 
    cp_elements(2210) <= OrReduce(cp_elements(2191) & cp_elements(2209));
    -- CP-element group 2211 fork  transition  bypass 
    -- predecessors 2210 
    -- successors 2212 2213 
    -- members (1) 
      -- 	branch_block_stmt_2042/merge_stmt_3435_PhiAck/$entry
      -- 
    cp_elements(2211) <= cp_elements(2210);
    -- CP-element group 2212 transition  input  bypass 
    -- predecessors 2211 
    -- successors 2214 
    -- members (1) 
      -- 	branch_block_stmt_2042/merge_stmt_3435_PhiAck/phi_stmt_3436_ack
      -- 
    phi_stmt_3436_ack_19078_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_3436_ack_0, ack => cp_elements(2212)); -- 
    -- CP-element group 2213 transition  input  bypass 
    -- predecessors 2211 
    -- successors 2214 
    -- members (1) 
      -- 	branch_block_stmt_2042/merge_stmt_3435_PhiAck/phi_stmt_3443_ack
      -- 
    phi_stmt_3443_ack_19079_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_3443_ack_0, ack => cp_elements(2213)); -- 
    -- CP-element group 2214 join  transition  bypass 
    -- predecessors 2212 2213 
    -- successors 56 
    -- members (1) 
      -- 	branch_block_stmt_2042/merge_stmt_3435_PhiAck/$exit
      -- 
    cp_element_group_2214: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_2214"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(2212) & cp_elements(2213);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(2214), clk => clk, reset => reset); --
    end block;
    -- CP-element group 2215 fork  transition  bypass 
    -- predecessors 950 
    -- successors 2216 2222 
    -- members (1) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi_udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi_PhiReq/$entry
      -- 
    cp_elements(2215) <= cp_elements(950);
    -- CP-element group 2216 fork  transition  bypass 
    -- predecessors 2215 
    -- successors 2217 2219 
    -- members (4) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi_udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi_PhiReq/phi_stmt_3498/$entry
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi_udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi_PhiReq/phi_stmt_3498/phi_stmt_3498_sources/$entry
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi_udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi_PhiReq/phi_stmt_3498/phi_stmt_3498_sources/type_cast_3501/$entry
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi_udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi_PhiReq/phi_stmt_3498/phi_stmt_3498_sources/type_cast_3501/SplitProtocol/$entry
      -- 
    cp_elements(2216) <= cp_elements(2215);
    -- CP-element group 2217 transition  output  bypass 
    -- predecessors 2216 
    -- successors 2218 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi_udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi_PhiReq/phi_stmt_3498/phi_stmt_3498_sources/type_cast_3501/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi_udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi_PhiReq/phi_stmt_3498/phi_stmt_3498_sources/type_cast_3501/SplitProtocol/Sample/rr
      -- 
    cp_elements(2217) <= cp_elements(2216);
    rr_19102_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2217), ack => type_cast_3501_inst_req_0); -- 
    -- CP-element group 2218 transition  input  bypass 
    -- predecessors 2217 
    -- successors 2221 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi_udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi_PhiReq/phi_stmt_3498/phi_stmt_3498_sources/type_cast_3501/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi_udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi_PhiReq/phi_stmt_3498/phi_stmt_3498_sources/type_cast_3501/SplitProtocol/Sample/ra
      -- 
    ra_19103_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3501_inst_ack_0, ack => cp_elements(2218)); -- 
    -- CP-element group 2219 transition  output  bypass 
    -- predecessors 2216 
    -- successors 2220 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi_udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi_PhiReq/phi_stmt_3498/phi_stmt_3498_sources/type_cast_3501/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi_udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi_PhiReq/phi_stmt_3498/phi_stmt_3498_sources/type_cast_3501/SplitProtocol/Update/cr
      -- 
    cp_elements(2219) <= cp_elements(2216);
    cr_19107_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2219), ack => type_cast_3501_inst_req_1); -- 
    -- CP-element group 2220 transition  input  bypass 
    -- predecessors 2219 
    -- successors 2221 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi_udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi_PhiReq/phi_stmt_3498/phi_stmt_3498_sources/type_cast_3501/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi_udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi_PhiReq/phi_stmt_3498/phi_stmt_3498_sources/type_cast_3501/SplitProtocol/Update/ca
      -- 
    ca_19108_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3501_inst_ack_1, ack => cp_elements(2220)); -- 
    -- CP-element group 2221 join  transition  output  bypass 
    -- predecessors 2218 2220 
    -- successors 2228 
    -- members (5) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi_udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi_PhiReq/phi_stmt_3498/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi_udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi_PhiReq/phi_stmt_3498/phi_stmt_3498_sources/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi_udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi_PhiReq/phi_stmt_3498/phi_stmt_3498_sources/type_cast_3501/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi_udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi_PhiReq/phi_stmt_3498/phi_stmt_3498_sources/type_cast_3501/SplitProtocol/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi_udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi_PhiReq/phi_stmt_3498/phi_stmt_3498_req
      -- 
    cp_element_group_2221: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_2221"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(2218) & cp_elements(2220);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(2221), clk => clk, reset => reset); --
    end block;
    phi_stmt_3498_req_19109_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2221), ack => phi_stmt_3498_req_0); -- 
    -- CP-element group 2222 fork  transition  bypass 
    -- predecessors 2215 
    -- successors 2223 2225 
    -- members (4) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi_udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi_PhiReq/phi_stmt_3494/$entry
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi_udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi_PhiReq/phi_stmt_3494/phi_stmt_3494_sources/$entry
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi_udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi_PhiReq/phi_stmt_3494/phi_stmt_3494_sources/type_cast_3497/$entry
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi_udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi_PhiReq/phi_stmt_3494/phi_stmt_3494_sources/type_cast_3497/SplitProtocol/$entry
      -- 
    cp_elements(2222) <= cp_elements(2215);
    -- CP-element group 2223 transition  output  bypass 
    -- predecessors 2222 
    -- successors 2224 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi_udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi_PhiReq/phi_stmt_3494/phi_stmt_3494_sources/type_cast_3497/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi_udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi_PhiReq/phi_stmt_3494/phi_stmt_3494_sources/type_cast_3497/SplitProtocol/Sample/rr
      -- 
    cp_elements(2223) <= cp_elements(2222);
    rr_19125_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2223), ack => type_cast_3497_inst_req_0); -- 
    -- CP-element group 2224 transition  input  bypass 
    -- predecessors 2223 
    -- successors 2227 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi_udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi_PhiReq/phi_stmt_3494/phi_stmt_3494_sources/type_cast_3497/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi_udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi_PhiReq/phi_stmt_3494/phi_stmt_3494_sources/type_cast_3497/SplitProtocol/Sample/ra
      -- 
    ra_19126_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3497_inst_ack_0, ack => cp_elements(2224)); -- 
    -- CP-element group 2225 transition  output  bypass 
    -- predecessors 2222 
    -- successors 2226 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi_udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi_PhiReq/phi_stmt_3494/phi_stmt_3494_sources/type_cast_3497/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi_udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi_PhiReq/phi_stmt_3494/phi_stmt_3494_sources/type_cast_3497/SplitProtocol/Update/cr
      -- 
    cp_elements(2225) <= cp_elements(2222);
    cr_19130_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2225), ack => type_cast_3497_inst_req_1); -- 
    -- CP-element group 2226 transition  input  bypass 
    -- predecessors 2225 
    -- successors 2227 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi_udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi_PhiReq/phi_stmt_3494/phi_stmt_3494_sources/type_cast_3497/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi_udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi_PhiReq/phi_stmt_3494/phi_stmt_3494_sources/type_cast_3497/SplitProtocol/Update/ca
      -- 
    ca_19131_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3497_inst_ack_1, ack => cp_elements(2226)); -- 
    -- CP-element group 2227 join  transition  output  bypass 
    -- predecessors 2224 2226 
    -- successors 2228 
    -- members (5) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi_udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi_PhiReq/phi_stmt_3494/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi_udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi_PhiReq/phi_stmt_3494/phi_stmt_3494_sources/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi_udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi_PhiReq/phi_stmt_3494/phi_stmt_3494_sources/type_cast_3497/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi_udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi_PhiReq/phi_stmt_3494/phi_stmt_3494_sources/type_cast_3497/SplitProtocol/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi_udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi_PhiReq/phi_stmt_3494/phi_stmt_3494_req
      -- 
    cp_element_group_2227: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_2227"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(2224) & cp_elements(2226);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(2227), clk => clk, reset => reset); --
    end block;
    phi_stmt_3494_req_19132_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2227), ack => phi_stmt_3494_req_0); -- 
    -- CP-element group 2228 join  transition  bypass 
    -- predecessors 2221 2227 
    -- successors 2229 
    -- members (1) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xi_udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi_PhiReq/$exit
      -- 
    cp_element_group_2228: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_2228"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(2221) & cp_elements(2227);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(2228), clk => clk, reset => reset); --
    end block;
    -- CP-element group 2229 place  bypass 
    -- predecessors 2228 
    -- successors 2230 
    -- members (1) 
      -- 	branch_block_stmt_2042/merge_stmt_3493_PhiReqMerge
      -- 
    cp_elements(2229) <= cp_elements(2228);
    -- CP-element group 2230 fork  transition  bypass 
    -- predecessors 2229 
    -- successors 2231 2232 
    -- members (1) 
      -- 	branch_block_stmt_2042/merge_stmt_3493_PhiAck/$entry
      -- 
    cp_elements(2230) <= cp_elements(2229);
    -- CP-element group 2231 transition  input  bypass 
    -- predecessors 2230 
    -- successors 2233 
    -- members (1) 
      -- 	branch_block_stmt_2042/merge_stmt_3493_PhiAck/phi_stmt_3494_ack
      -- 
    phi_stmt_3494_ack_19137_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_3494_ack_0, ack => cp_elements(2231)); -- 
    -- CP-element group 2232 transition  input  bypass 
    -- predecessors 2230 
    -- successors 2233 
    -- members (1) 
      -- 	branch_block_stmt_2042/merge_stmt_3493_PhiAck/phi_stmt_3498_ack
      -- 
    phi_stmt_3498_ack_19138_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_3498_ack_0, ack => cp_elements(2232)); -- 
    -- CP-element group 2233 join  transition  bypass 
    -- predecessors 2231 2232 
    -- successors 58 
    -- members (1) 
      -- 	branch_block_stmt_2042/merge_stmt_3493_PhiAck/$exit
      -- 
    cp_element_group_2233: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_2233"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(2231) & cp_elements(2232);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(2233), clk => clk, reset => reset); --
    end block;
    -- CP-element group 2234 fork  transition  bypass 
    -- predecessors 916 
    -- successors 2235 2247 
    -- members (1) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xpreheaderx_xix_xi_xx_xcritedgex_xix_xi_PhiReq/$entry
      -- 
    cp_elements(2234) <= cp_elements(916);
    -- CP-element group 2235 fork  transition  bypass 
    -- predecessors 2234 
    -- successors 2236 2240 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xpreheaderx_xix_xi_xx_xcritedgex_xix_xi_PhiReq/phi_stmt_3521/$entry
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xpreheaderx_xix_xi_xx_xcritedgex_xix_xi_PhiReq/phi_stmt_3521/phi_stmt_3521_sources/$entry
      -- 
    cp_elements(2235) <= cp_elements(2234);
    -- CP-element group 2236 fork  transition  bypass 
    -- predecessors 2235 
    -- successors 2237 2238 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xpreheaderx_xix_xi_xx_xcritedgex_xix_xi_PhiReq/phi_stmt_3521/phi_stmt_3521_sources/type_cast_3524/$entry
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xpreheaderx_xix_xi_xx_xcritedgex_xix_xi_PhiReq/phi_stmt_3521/phi_stmt_3521_sources/type_cast_3524/SplitProtocol/$entry
      -- 
    cp_elements(2236) <= cp_elements(2235);
    -- CP-element group 2237 transition  bypass 
    -- predecessors 2236 
    -- successors 2239 
    -- members (4) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xpreheaderx_xix_xi_xx_xcritedgex_xix_xi_PhiReq/phi_stmt_3521/phi_stmt_3521_sources/type_cast_3524/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xpreheaderx_xix_xi_xx_xcritedgex_xix_xi_PhiReq/phi_stmt_3521/phi_stmt_3521_sources/type_cast_3524/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xpreheaderx_xix_xi_xx_xcritedgex_xix_xi_PhiReq/phi_stmt_3521/phi_stmt_3521_sources/type_cast_3524/SplitProtocol/Sample/rr
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xpreheaderx_xix_xi_xx_xcritedgex_xix_xi_PhiReq/phi_stmt_3521/phi_stmt_3521_sources/type_cast_3524/SplitProtocol/Sample/ra
      -- 
    cp_elements(2237) <= cp_elements(2236);
    -- CP-element group 2238 transition  bypass 
    -- predecessors 2236 
    -- successors 2239 
    -- members (4) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xpreheaderx_xix_xi_xx_xcritedgex_xix_xi_PhiReq/phi_stmt_3521/phi_stmt_3521_sources/type_cast_3524/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xpreheaderx_xix_xi_xx_xcritedgex_xix_xi_PhiReq/phi_stmt_3521/phi_stmt_3521_sources/type_cast_3524/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xpreheaderx_xix_xi_xx_xcritedgex_xix_xi_PhiReq/phi_stmt_3521/phi_stmt_3521_sources/type_cast_3524/SplitProtocol/Update/cr
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xpreheaderx_xix_xi_xx_xcritedgex_xix_xi_PhiReq/phi_stmt_3521/phi_stmt_3521_sources/type_cast_3524/SplitProtocol/Update/ca
      -- 
    cp_elements(2238) <= cp_elements(2236);
    -- CP-element group 2239 join  transition  bypass 
    -- predecessors 2237 2238 
    -- successors 2246 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xpreheaderx_xix_xi_xx_xcritedgex_xix_xi_PhiReq/phi_stmt_3521/phi_stmt_3521_sources/type_cast_3524/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xpreheaderx_xix_xi_xx_xcritedgex_xix_xi_PhiReq/phi_stmt_3521/phi_stmt_3521_sources/type_cast_3524/SplitProtocol/$exit
      -- 
    cp_element_group_2239: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_2239"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(2237) & cp_elements(2238);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(2239), clk => clk, reset => reset); --
    end block;
    -- CP-element group 2240 fork  transition  bypass 
    -- predecessors 2235 
    -- successors 2241 2243 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xpreheaderx_xix_xi_xx_xcritedgex_xix_xi_PhiReq/phi_stmt_3521/phi_stmt_3521_sources/type_cast_3526/$entry
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xpreheaderx_xix_xi_xx_xcritedgex_xix_xi_PhiReq/phi_stmt_3521/phi_stmt_3521_sources/type_cast_3526/SplitProtocol/$entry
      -- 
    cp_elements(2240) <= cp_elements(2235);
    -- CP-element group 2241 transition  output  bypass 
    -- predecessors 2240 
    -- successors 2242 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xpreheaderx_xix_xi_xx_xcritedgex_xix_xi_PhiReq/phi_stmt_3521/phi_stmt_3521_sources/type_cast_3526/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xpreheaderx_xix_xi_xx_xcritedgex_xix_xi_PhiReq/phi_stmt_3521/phi_stmt_3521_sources/type_cast_3526/SplitProtocol/Sample/rr
      -- 
    cp_elements(2241) <= cp_elements(2240);
    rr_19173_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2241), ack => type_cast_3526_inst_req_0); -- 
    -- CP-element group 2242 transition  input  bypass 
    -- predecessors 2241 
    -- successors 2245 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xpreheaderx_xix_xi_xx_xcritedgex_xix_xi_PhiReq/phi_stmt_3521/phi_stmt_3521_sources/type_cast_3526/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xpreheaderx_xix_xi_xx_xcritedgex_xix_xi_PhiReq/phi_stmt_3521/phi_stmt_3521_sources/type_cast_3526/SplitProtocol/Sample/ra
      -- 
    ra_19174_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3526_inst_ack_0, ack => cp_elements(2242)); -- 
    -- CP-element group 2243 transition  output  bypass 
    -- predecessors 2240 
    -- successors 2244 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xpreheaderx_xix_xi_xx_xcritedgex_xix_xi_PhiReq/phi_stmt_3521/phi_stmt_3521_sources/type_cast_3526/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xpreheaderx_xix_xi_xx_xcritedgex_xix_xi_PhiReq/phi_stmt_3521/phi_stmt_3521_sources/type_cast_3526/SplitProtocol/Update/cr
      -- 
    cp_elements(2243) <= cp_elements(2240);
    cr_19178_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2243), ack => type_cast_3526_inst_req_1); -- 
    -- CP-element group 2244 transition  input  bypass 
    -- predecessors 2243 
    -- successors 2245 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xpreheaderx_xix_xi_xx_xcritedgex_xix_xi_PhiReq/phi_stmt_3521/phi_stmt_3521_sources/type_cast_3526/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xpreheaderx_xix_xi_xx_xcritedgex_xix_xi_PhiReq/phi_stmt_3521/phi_stmt_3521_sources/type_cast_3526/SplitProtocol/Update/ca
      -- 
    ca_19179_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3526_inst_ack_1, ack => cp_elements(2244)); -- 
    -- CP-element group 2245 join  transition  bypass 
    -- predecessors 2242 2244 
    -- successors 2246 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xpreheaderx_xix_xi_xx_xcritedgex_xix_xi_PhiReq/phi_stmt_3521/phi_stmt_3521_sources/type_cast_3526/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xpreheaderx_xix_xi_xx_xcritedgex_xix_xi_PhiReq/phi_stmt_3521/phi_stmt_3521_sources/type_cast_3526/SplitProtocol/$exit
      -- 
    cp_element_group_2245: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_2245"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(2242) & cp_elements(2244);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(2245), clk => clk, reset => reset); --
    end block;
    -- CP-element group 2246 join  transition  output  bypass 
    -- predecessors 2239 2245 
    -- successors 2259 
    -- members (3) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xpreheaderx_xix_xi_xx_xcritedgex_xix_xi_PhiReq/phi_stmt_3521/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xpreheaderx_xix_xi_xx_xcritedgex_xix_xi_PhiReq/phi_stmt_3521/phi_stmt_3521_sources/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xpreheaderx_xix_xi_xx_xcritedgex_xix_xi_PhiReq/phi_stmt_3521/phi_stmt_3521_req
      -- 
    cp_element_group_2246: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_2246"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(2239) & cp_elements(2245);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(2246), clk => clk, reset => reset); --
    end block;
    phi_stmt_3521_req_19180_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2246), ack => phi_stmt_3521_req_1); -- 
    -- CP-element group 2247 fork  transition  bypass 
    -- predecessors 2234 
    -- successors 2248 2252 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xpreheaderx_xix_xi_xx_xcritedgex_xix_xi_PhiReq/phi_stmt_3527/$entry
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xpreheaderx_xix_xi_xx_xcritedgex_xix_xi_PhiReq/phi_stmt_3527/phi_stmt_3527_sources/$entry
      -- 
    cp_elements(2247) <= cp_elements(2234);
    -- CP-element group 2248 fork  transition  bypass 
    -- predecessors 2247 
    -- successors 2249 2250 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xpreheaderx_xix_xi_xx_xcritedgex_xix_xi_PhiReq/phi_stmt_3527/phi_stmt_3527_sources/type_cast_3530/$entry
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xpreheaderx_xix_xi_xx_xcritedgex_xix_xi_PhiReq/phi_stmt_3527/phi_stmt_3527_sources/type_cast_3530/SplitProtocol/$entry
      -- 
    cp_elements(2248) <= cp_elements(2247);
    -- CP-element group 2249 transition  bypass 
    -- predecessors 2248 
    -- successors 2251 
    -- members (4) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xpreheaderx_xix_xi_xx_xcritedgex_xix_xi_PhiReq/phi_stmt_3527/phi_stmt_3527_sources/type_cast_3530/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xpreheaderx_xix_xi_xx_xcritedgex_xix_xi_PhiReq/phi_stmt_3527/phi_stmt_3527_sources/type_cast_3530/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xpreheaderx_xix_xi_xx_xcritedgex_xix_xi_PhiReq/phi_stmt_3527/phi_stmt_3527_sources/type_cast_3530/SplitProtocol/Sample/rr
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xpreheaderx_xix_xi_xx_xcritedgex_xix_xi_PhiReq/phi_stmt_3527/phi_stmt_3527_sources/type_cast_3530/SplitProtocol/Sample/ra
      -- 
    cp_elements(2249) <= cp_elements(2248);
    -- CP-element group 2250 transition  bypass 
    -- predecessors 2248 
    -- successors 2251 
    -- members (4) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xpreheaderx_xix_xi_xx_xcritedgex_xix_xi_PhiReq/phi_stmt_3527/phi_stmt_3527_sources/type_cast_3530/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xpreheaderx_xix_xi_xx_xcritedgex_xix_xi_PhiReq/phi_stmt_3527/phi_stmt_3527_sources/type_cast_3530/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xpreheaderx_xix_xi_xx_xcritedgex_xix_xi_PhiReq/phi_stmt_3527/phi_stmt_3527_sources/type_cast_3530/SplitProtocol/Update/cr
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xpreheaderx_xix_xi_xx_xcritedgex_xix_xi_PhiReq/phi_stmt_3527/phi_stmt_3527_sources/type_cast_3530/SplitProtocol/Update/ca
      -- 
    cp_elements(2250) <= cp_elements(2248);
    -- CP-element group 2251 join  transition  bypass 
    -- predecessors 2249 2250 
    -- successors 2258 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xpreheaderx_xix_xi_xx_xcritedgex_xix_xi_PhiReq/phi_stmt_3527/phi_stmt_3527_sources/type_cast_3530/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xpreheaderx_xix_xi_xx_xcritedgex_xix_xi_PhiReq/phi_stmt_3527/phi_stmt_3527_sources/type_cast_3530/SplitProtocol/$exit
      -- 
    cp_element_group_2251: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_2251"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(2249) & cp_elements(2250);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(2251), clk => clk, reset => reset); --
    end block;
    -- CP-element group 2252 fork  transition  bypass 
    -- predecessors 2247 
    -- successors 2253 2255 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xpreheaderx_xix_xi_xx_xcritedgex_xix_xi_PhiReq/phi_stmt_3527/phi_stmt_3527_sources/type_cast_3532/$entry
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xpreheaderx_xix_xi_xx_xcritedgex_xix_xi_PhiReq/phi_stmt_3527/phi_stmt_3527_sources/type_cast_3532/SplitProtocol/$entry
      -- 
    cp_elements(2252) <= cp_elements(2247);
    -- CP-element group 2253 transition  output  bypass 
    -- predecessors 2252 
    -- successors 2254 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xpreheaderx_xix_xi_xx_xcritedgex_xix_xi_PhiReq/phi_stmt_3527/phi_stmt_3527_sources/type_cast_3532/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xpreheaderx_xix_xi_xx_xcritedgex_xix_xi_PhiReq/phi_stmt_3527/phi_stmt_3527_sources/type_cast_3532/SplitProtocol/Sample/rr
      -- 
    cp_elements(2253) <= cp_elements(2252);
    rr_19212_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2253), ack => type_cast_3532_inst_req_0); -- 
    -- CP-element group 2254 transition  input  bypass 
    -- predecessors 2253 
    -- successors 2257 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xpreheaderx_xix_xi_xx_xcritedgex_xix_xi_PhiReq/phi_stmt_3527/phi_stmt_3527_sources/type_cast_3532/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xpreheaderx_xix_xi_xx_xcritedgex_xix_xi_PhiReq/phi_stmt_3527/phi_stmt_3527_sources/type_cast_3532/SplitProtocol/Sample/ra
      -- 
    ra_19213_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3532_inst_ack_0, ack => cp_elements(2254)); -- 
    -- CP-element group 2255 transition  output  bypass 
    -- predecessors 2252 
    -- successors 2256 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xpreheaderx_xix_xi_xx_xcritedgex_xix_xi_PhiReq/phi_stmt_3527/phi_stmt_3527_sources/type_cast_3532/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xpreheaderx_xix_xi_xx_xcritedgex_xix_xi_PhiReq/phi_stmt_3527/phi_stmt_3527_sources/type_cast_3532/SplitProtocol/Update/cr
      -- 
    cp_elements(2255) <= cp_elements(2252);
    cr_19217_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2255), ack => type_cast_3532_inst_req_1); -- 
    -- CP-element group 2256 transition  input  bypass 
    -- predecessors 2255 
    -- successors 2257 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xpreheaderx_xix_xi_xx_xcritedgex_xix_xi_PhiReq/phi_stmt_3527/phi_stmt_3527_sources/type_cast_3532/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xpreheaderx_xix_xi_xx_xcritedgex_xix_xi_PhiReq/phi_stmt_3527/phi_stmt_3527_sources/type_cast_3532/SplitProtocol/Update/ca
      -- 
    ca_19218_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3532_inst_ack_1, ack => cp_elements(2256)); -- 
    -- CP-element group 2257 join  transition  bypass 
    -- predecessors 2254 2256 
    -- successors 2258 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xpreheaderx_xix_xi_xx_xcritedgex_xix_xi_PhiReq/phi_stmt_3527/phi_stmt_3527_sources/type_cast_3532/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xpreheaderx_xix_xi_xx_xcritedgex_xix_xi_PhiReq/phi_stmt_3527/phi_stmt_3527_sources/type_cast_3532/SplitProtocol/$exit
      -- 
    cp_element_group_2257: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_2257"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(2254) & cp_elements(2256);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(2257), clk => clk, reset => reset); --
    end block;
    -- CP-element group 2258 join  transition  output  bypass 
    -- predecessors 2251 2257 
    -- successors 2259 
    -- members (3) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xpreheaderx_xix_xi_xx_xcritedgex_xix_xi_PhiReq/phi_stmt_3527/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xpreheaderx_xix_xi_xx_xcritedgex_xix_xi_PhiReq/phi_stmt_3527/phi_stmt_3527_sources/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xpreheaderx_xix_xi_xx_xcritedgex_xix_xi_PhiReq/phi_stmt_3527/phi_stmt_3527_req
      -- 
    cp_element_group_2258: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_2258"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(2251) & cp_elements(2257);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(2258), clk => clk, reset => reset); --
    end block;
    phi_stmt_3527_req_19219_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2258), ack => phi_stmt_3527_req_1); -- 
    -- CP-element group 2259 join  transition  bypass 
    -- predecessors 2246 2258 
    -- successors 2286 
    -- members (1) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xpreheaderx_xix_xi_xx_xcritedgex_xix_xi_PhiReq/$exit
      -- 
    cp_element_group_2259: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_2259"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(2246) & cp_elements(2258);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(2259), clk => clk, reset => reset); --
    end block;
    -- CP-element group 2260 fork  transition  bypass 
    -- predecessors 965 
    -- successors 2261 2273 
    -- members (1) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi_xx_xcritedgex_xix_xi_PhiReq/$entry
      -- 
    cp_elements(2260) <= cp_elements(965);
    -- CP-element group 2261 fork  transition  bypass 
    -- predecessors 2260 
    -- successors 2262 2268 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi_xx_xcritedgex_xix_xi_PhiReq/phi_stmt_3521/$entry
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi_xx_xcritedgex_xix_xi_PhiReq/phi_stmt_3521/phi_stmt_3521_sources/$entry
      -- 
    cp_elements(2261) <= cp_elements(2260);
    -- CP-element group 2262 fork  transition  bypass 
    -- predecessors 2261 
    -- successors 2263 2265 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi_xx_xcritedgex_xix_xi_PhiReq/phi_stmt_3521/phi_stmt_3521_sources/type_cast_3524/$entry
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi_xx_xcritedgex_xix_xi_PhiReq/phi_stmt_3521/phi_stmt_3521_sources/type_cast_3524/SplitProtocol/$entry
      -- 
    cp_elements(2262) <= cp_elements(2261);
    -- CP-element group 2263 transition  output  bypass 
    -- predecessors 2262 
    -- successors 2264 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi_xx_xcritedgex_xix_xi_PhiReq/phi_stmt_3521/phi_stmt_3521_sources/type_cast_3524/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi_xx_xcritedgex_xix_xi_PhiReq/phi_stmt_3521/phi_stmt_3521_sources/type_cast_3524/SplitProtocol/Sample/rr
      -- 
    cp_elements(2263) <= cp_elements(2262);
    rr_19238_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2263), ack => type_cast_3524_inst_req_0); -- 
    -- CP-element group 2264 transition  input  bypass 
    -- predecessors 2263 
    -- successors 2267 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi_xx_xcritedgex_xix_xi_PhiReq/phi_stmt_3521/phi_stmt_3521_sources/type_cast_3524/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi_xx_xcritedgex_xix_xi_PhiReq/phi_stmt_3521/phi_stmt_3521_sources/type_cast_3524/SplitProtocol/Sample/ra
      -- 
    ra_19239_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3524_inst_ack_0, ack => cp_elements(2264)); -- 
    -- CP-element group 2265 transition  output  bypass 
    -- predecessors 2262 
    -- successors 2266 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi_xx_xcritedgex_xix_xi_PhiReq/phi_stmt_3521/phi_stmt_3521_sources/type_cast_3524/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi_xx_xcritedgex_xix_xi_PhiReq/phi_stmt_3521/phi_stmt_3521_sources/type_cast_3524/SplitProtocol/Update/cr
      -- 
    cp_elements(2265) <= cp_elements(2262);
    cr_19243_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2265), ack => type_cast_3524_inst_req_1); -- 
    -- CP-element group 2266 transition  input  bypass 
    -- predecessors 2265 
    -- successors 2267 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi_xx_xcritedgex_xix_xi_PhiReq/phi_stmt_3521/phi_stmt_3521_sources/type_cast_3524/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi_xx_xcritedgex_xix_xi_PhiReq/phi_stmt_3521/phi_stmt_3521_sources/type_cast_3524/SplitProtocol/Update/ca
      -- 
    ca_19244_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3524_inst_ack_1, ack => cp_elements(2266)); -- 
    -- CP-element group 2267 join  transition  bypass 
    -- predecessors 2264 2266 
    -- successors 2272 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi_xx_xcritedgex_xix_xi_PhiReq/phi_stmt_3521/phi_stmt_3521_sources/type_cast_3524/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi_xx_xcritedgex_xix_xi_PhiReq/phi_stmt_3521/phi_stmt_3521_sources/type_cast_3524/SplitProtocol/$exit
      -- 
    cp_element_group_2267: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_2267"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(2264) & cp_elements(2266);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(2267), clk => clk, reset => reset); --
    end block;
    -- CP-element group 2268 fork  transition  bypass 
    -- predecessors 2261 
    -- successors 2269 2270 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi_xx_xcritedgex_xix_xi_PhiReq/phi_stmt_3521/phi_stmt_3521_sources/type_cast_3526/$entry
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi_xx_xcritedgex_xix_xi_PhiReq/phi_stmt_3521/phi_stmt_3521_sources/type_cast_3526/SplitProtocol/$entry
      -- 
    cp_elements(2268) <= cp_elements(2261);
    -- CP-element group 2269 transition  bypass 
    -- predecessors 2268 
    -- successors 2271 
    -- members (4) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi_xx_xcritedgex_xix_xi_PhiReq/phi_stmt_3521/phi_stmt_3521_sources/type_cast_3526/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi_xx_xcritedgex_xix_xi_PhiReq/phi_stmt_3521/phi_stmt_3521_sources/type_cast_3526/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi_xx_xcritedgex_xix_xi_PhiReq/phi_stmt_3521/phi_stmt_3521_sources/type_cast_3526/SplitProtocol/Sample/rr
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi_xx_xcritedgex_xix_xi_PhiReq/phi_stmt_3521/phi_stmt_3521_sources/type_cast_3526/SplitProtocol/Sample/ra
      -- 
    cp_elements(2269) <= cp_elements(2268);
    -- CP-element group 2270 transition  bypass 
    -- predecessors 2268 
    -- successors 2271 
    -- members (4) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi_xx_xcritedgex_xix_xi_PhiReq/phi_stmt_3521/phi_stmt_3521_sources/type_cast_3526/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi_xx_xcritedgex_xix_xi_PhiReq/phi_stmt_3521/phi_stmt_3521_sources/type_cast_3526/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi_xx_xcritedgex_xix_xi_PhiReq/phi_stmt_3521/phi_stmt_3521_sources/type_cast_3526/SplitProtocol/Update/cr
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi_xx_xcritedgex_xix_xi_PhiReq/phi_stmt_3521/phi_stmt_3521_sources/type_cast_3526/SplitProtocol/Update/ca
      -- 
    cp_elements(2270) <= cp_elements(2268);
    -- CP-element group 2271 join  transition  bypass 
    -- predecessors 2269 2270 
    -- successors 2272 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi_xx_xcritedgex_xix_xi_PhiReq/phi_stmt_3521/phi_stmt_3521_sources/type_cast_3526/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi_xx_xcritedgex_xix_xi_PhiReq/phi_stmt_3521/phi_stmt_3521_sources/type_cast_3526/SplitProtocol/$exit
      -- 
    cp_element_group_2271: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_2271"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(2269) & cp_elements(2270);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(2271), clk => clk, reset => reset); --
    end block;
    -- CP-element group 2272 join  transition  output  bypass 
    -- predecessors 2267 2271 
    -- successors 2285 
    -- members (3) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi_xx_xcritedgex_xix_xi_PhiReq/phi_stmt_3521/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi_xx_xcritedgex_xix_xi_PhiReq/phi_stmt_3521/phi_stmt_3521_sources/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi_xx_xcritedgex_xix_xi_PhiReq/phi_stmt_3521/phi_stmt_3521_req
      -- 
    cp_element_group_2272: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_2272"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(2267) & cp_elements(2271);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(2272), clk => clk, reset => reset); --
    end block;
    phi_stmt_3521_req_19261_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2272), ack => phi_stmt_3521_req_0); -- 
    -- CP-element group 2273 fork  transition  bypass 
    -- predecessors 2260 
    -- successors 2274 2280 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi_xx_xcritedgex_xix_xi_PhiReq/phi_stmt_3527/$entry
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi_xx_xcritedgex_xix_xi_PhiReq/phi_stmt_3527/phi_stmt_3527_sources/$entry
      -- 
    cp_elements(2273) <= cp_elements(2260);
    -- CP-element group 2274 fork  transition  bypass 
    -- predecessors 2273 
    -- successors 2275 2277 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi_xx_xcritedgex_xix_xi_PhiReq/phi_stmt_3527/phi_stmt_3527_sources/type_cast_3530/$entry
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi_xx_xcritedgex_xix_xi_PhiReq/phi_stmt_3527/phi_stmt_3527_sources/type_cast_3530/SplitProtocol/$entry
      -- 
    cp_elements(2274) <= cp_elements(2273);
    -- CP-element group 2275 transition  output  bypass 
    -- predecessors 2274 
    -- successors 2276 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi_xx_xcritedgex_xix_xi_PhiReq/phi_stmt_3527/phi_stmt_3527_sources/type_cast_3530/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi_xx_xcritedgex_xix_xi_PhiReq/phi_stmt_3527/phi_stmt_3527_sources/type_cast_3530/SplitProtocol/Sample/rr
      -- 
    cp_elements(2275) <= cp_elements(2274);
    rr_19277_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2275), ack => type_cast_3530_inst_req_0); -- 
    -- CP-element group 2276 transition  input  bypass 
    -- predecessors 2275 
    -- successors 2279 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi_xx_xcritedgex_xix_xi_PhiReq/phi_stmt_3527/phi_stmt_3527_sources/type_cast_3530/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi_xx_xcritedgex_xix_xi_PhiReq/phi_stmt_3527/phi_stmt_3527_sources/type_cast_3530/SplitProtocol/Sample/ra
      -- 
    ra_19278_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3530_inst_ack_0, ack => cp_elements(2276)); -- 
    -- CP-element group 2277 transition  output  bypass 
    -- predecessors 2274 
    -- successors 2278 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi_xx_xcritedgex_xix_xi_PhiReq/phi_stmt_3527/phi_stmt_3527_sources/type_cast_3530/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi_xx_xcritedgex_xix_xi_PhiReq/phi_stmt_3527/phi_stmt_3527_sources/type_cast_3530/SplitProtocol/Update/cr
      -- 
    cp_elements(2277) <= cp_elements(2274);
    cr_19282_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2277), ack => type_cast_3530_inst_req_1); -- 
    -- CP-element group 2278 transition  input  bypass 
    -- predecessors 2277 
    -- successors 2279 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi_xx_xcritedgex_xix_xi_PhiReq/phi_stmt_3527/phi_stmt_3527_sources/type_cast_3530/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi_xx_xcritedgex_xix_xi_PhiReq/phi_stmt_3527/phi_stmt_3527_sources/type_cast_3530/SplitProtocol/Update/ca
      -- 
    ca_19283_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3530_inst_ack_1, ack => cp_elements(2278)); -- 
    -- CP-element group 2279 join  transition  bypass 
    -- predecessors 2276 2278 
    -- successors 2284 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi_xx_xcritedgex_xix_xi_PhiReq/phi_stmt_3527/phi_stmt_3527_sources/type_cast_3530/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi_xx_xcritedgex_xix_xi_PhiReq/phi_stmt_3527/phi_stmt_3527_sources/type_cast_3530/SplitProtocol/$exit
      -- 
    cp_element_group_2279: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_2279"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(2276) & cp_elements(2278);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(2279), clk => clk, reset => reset); --
    end block;
    -- CP-element group 2280 fork  transition  bypass 
    -- predecessors 2273 
    -- successors 2281 2282 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi_xx_xcritedgex_xix_xi_PhiReq/phi_stmt_3527/phi_stmt_3527_sources/type_cast_3532/$entry
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi_xx_xcritedgex_xix_xi_PhiReq/phi_stmt_3527/phi_stmt_3527_sources/type_cast_3532/SplitProtocol/$entry
      -- 
    cp_elements(2280) <= cp_elements(2273);
    -- CP-element group 2281 transition  bypass 
    -- predecessors 2280 
    -- successors 2283 
    -- members (4) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi_xx_xcritedgex_xix_xi_PhiReq/phi_stmt_3527/phi_stmt_3527_sources/type_cast_3532/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi_xx_xcritedgex_xix_xi_PhiReq/phi_stmt_3527/phi_stmt_3527_sources/type_cast_3532/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi_xx_xcritedgex_xix_xi_PhiReq/phi_stmt_3527/phi_stmt_3527_sources/type_cast_3532/SplitProtocol/Sample/rr
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi_xx_xcritedgex_xix_xi_PhiReq/phi_stmt_3527/phi_stmt_3527_sources/type_cast_3532/SplitProtocol/Sample/ra
      -- 
    cp_elements(2281) <= cp_elements(2280);
    -- CP-element group 2282 transition  bypass 
    -- predecessors 2280 
    -- successors 2283 
    -- members (4) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi_xx_xcritedgex_xix_xi_PhiReq/phi_stmt_3527/phi_stmt_3527_sources/type_cast_3532/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi_xx_xcritedgex_xix_xi_PhiReq/phi_stmt_3527/phi_stmt_3527_sources/type_cast_3532/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi_xx_xcritedgex_xix_xi_PhiReq/phi_stmt_3527/phi_stmt_3527_sources/type_cast_3532/SplitProtocol/Update/cr
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi_xx_xcritedgex_xix_xi_PhiReq/phi_stmt_3527/phi_stmt_3527_sources/type_cast_3532/SplitProtocol/Update/ca
      -- 
    cp_elements(2282) <= cp_elements(2280);
    -- CP-element group 2283 join  transition  bypass 
    -- predecessors 2281 2282 
    -- successors 2284 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi_xx_xcritedgex_xix_xi_PhiReq/phi_stmt_3527/phi_stmt_3527_sources/type_cast_3532/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi_xx_xcritedgex_xix_xi_PhiReq/phi_stmt_3527/phi_stmt_3527_sources/type_cast_3532/SplitProtocol/$exit
      -- 
    cp_element_group_2283: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_2283"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(2281) & cp_elements(2282);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(2283), clk => clk, reset => reset); --
    end block;
    -- CP-element group 2284 join  transition  output  bypass 
    -- predecessors 2279 2283 
    -- successors 2285 
    -- members (3) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi_xx_xcritedgex_xix_xi_PhiReq/phi_stmt_3527/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi_xx_xcritedgex_xix_xi_PhiReq/phi_stmt_3527/phi_stmt_3527_sources/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi_xx_xcritedgex_xix_xi_PhiReq/phi_stmt_3527/phi_stmt_3527_req
      -- 
    cp_element_group_2284: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_2284"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(2279) & cp_elements(2283);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(2284), clk => clk, reset => reset); --
    end block;
    phi_stmt_3527_req_19300_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2284), ack => phi_stmt_3527_req_0); -- 
    -- CP-element group 2285 join  transition  bypass 
    -- predecessors 2272 2284 
    -- successors 2286 
    -- members (1) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi_xx_xcritedgex_xix_xi_PhiReq/$exit
      -- 
    cp_element_group_2285: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_2285"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(2272) & cp_elements(2284);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(2285), clk => clk, reset => reset); --
    end block;
    -- CP-element group 2286 merge  place  bypass 
    -- predecessors 2259 2285 
    -- successors 2287 
    -- members (1) 
      -- 	branch_block_stmt_2042/merge_stmt_3520_PhiReqMerge
      -- 
    cp_elements(2286) <= OrReduce(cp_elements(2259) & cp_elements(2285));
    -- CP-element group 2287 fork  transition  bypass 
    -- predecessors 2286 
    -- successors 2288 2289 
    -- members (1) 
      -- 	branch_block_stmt_2042/merge_stmt_3520_PhiAck/$entry
      -- 
    cp_elements(2287) <= cp_elements(2286);
    -- CP-element group 2288 transition  input  bypass 
    -- predecessors 2287 
    -- successors 2290 
    -- members (1) 
      -- 	branch_block_stmt_2042/merge_stmt_3520_PhiAck/phi_stmt_3521_ack
      -- 
    phi_stmt_3521_ack_19305_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_3521_ack_0, ack => cp_elements(2288)); -- 
    -- CP-element group 2289 transition  input  bypass 
    -- predecessors 2287 
    -- successors 2290 
    -- members (1) 
      -- 	branch_block_stmt_2042/merge_stmt_3520_PhiAck/phi_stmt_3527_ack
      -- 
    phi_stmt_3527_ack_19306_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_3527_ack_0, ack => cp_elements(2289)); -- 
    -- CP-element group 2290 join  transition  bypass 
    -- predecessors 2288 2289 
    -- successors 59 
    -- members (1) 
      -- 	branch_block_stmt_2042/merge_stmt_3520_PhiAck/$exit
      -- 
    cp_element_group_2290: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_2290"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(2288) & cp_elements(2289);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(2290), clk => clk, reset => reset); --
    end block;
    -- CP-element group 2291 transition  bypass 
    -- predecessors 752 
    -- successors 2293 
    -- members (4) 
      -- 	branch_block_stmt_2042/omega_calcx_xexit_iq_err_calcx_xexit_PhiReq/phi_stmt_3568/phi_stmt_3568_sources/type_cast_3571/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_2042/omega_calcx_xexit_iq_err_calcx_xexit_PhiReq/phi_stmt_3568/phi_stmt_3568_sources/type_cast_3571/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_2042/omega_calcx_xexit_iq_err_calcx_xexit_PhiReq/phi_stmt_3568/phi_stmt_3568_sources/type_cast_3571/SplitProtocol/Sample/rr
      -- 	branch_block_stmt_2042/omega_calcx_xexit_iq_err_calcx_xexit_PhiReq/phi_stmt_3568/phi_stmt_3568_sources/type_cast_3571/SplitProtocol/Sample/ra
      -- 
    cp_elements(2291) <= cp_elements(752);
    -- CP-element group 2292 transition  bypass 
    -- predecessors 752 
    -- successors 2293 
    -- members (4) 
      -- 	branch_block_stmt_2042/omega_calcx_xexit_iq_err_calcx_xexit_PhiReq/phi_stmt_3568/phi_stmt_3568_sources/type_cast_3571/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_2042/omega_calcx_xexit_iq_err_calcx_xexit_PhiReq/phi_stmt_3568/phi_stmt_3568_sources/type_cast_3571/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_2042/omega_calcx_xexit_iq_err_calcx_xexit_PhiReq/phi_stmt_3568/phi_stmt_3568_sources/type_cast_3571/SplitProtocol/Update/cr
      -- 	branch_block_stmt_2042/omega_calcx_xexit_iq_err_calcx_xexit_PhiReq/phi_stmt_3568/phi_stmt_3568_sources/type_cast_3571/SplitProtocol/Update/ca
      -- 
    cp_elements(2292) <= cp_elements(752);
    -- CP-element group 2293 join  transition  output  bypass 
    -- predecessors 2291 2292 
    -- successors 2299 
    -- members (6) 
      -- 	branch_block_stmt_2042/omega_calcx_xexit_iq_err_calcx_xexit_PhiReq/$exit
      -- 	branch_block_stmt_2042/omega_calcx_xexit_iq_err_calcx_xexit_PhiReq/phi_stmt_3568/$exit
      -- 	branch_block_stmt_2042/omega_calcx_xexit_iq_err_calcx_xexit_PhiReq/phi_stmt_3568/phi_stmt_3568_sources/$exit
      -- 	branch_block_stmt_2042/omega_calcx_xexit_iq_err_calcx_xexit_PhiReq/phi_stmt_3568/phi_stmt_3568_sources/type_cast_3571/$exit
      -- 	branch_block_stmt_2042/omega_calcx_xexit_iq_err_calcx_xexit_PhiReq/phi_stmt_3568/phi_stmt_3568_sources/type_cast_3571/SplitProtocol/$exit
      -- 	branch_block_stmt_2042/omega_calcx_xexit_iq_err_calcx_xexit_PhiReq/phi_stmt_3568/phi_stmt_3568_req
      -- 
    cp_element_group_2293: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_2293"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(2291) & cp_elements(2292);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(2293), clk => clk, reset => reset); --
    end block;
    phi_stmt_3568_req_19332_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2293), ack => phi_stmt_3568_req_1); -- 
    -- CP-element group 2294 transition  output  bypass 
    -- predecessors 989 
    -- successors 2295 
    -- members (2) 
      -- 	branch_block_stmt_2042/xx_xcritedgex_xix_xi_iq_err_calcx_xexit_PhiReq/phi_stmt_3568/phi_stmt_3568_sources/type_cast_3571/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_2042/xx_xcritedgex_xix_xi_iq_err_calcx_xexit_PhiReq/phi_stmt_3568/phi_stmt_3568_sources/type_cast_3571/SplitProtocol/Sample/rr
      -- 
    cp_elements(2294) <= cp_elements(989);
    rr_19351_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2294), ack => type_cast_3571_inst_req_0); -- 
    -- CP-element group 2295 transition  input  bypass 
    -- predecessors 2294 
    -- successors 2298 
    -- members (2) 
      -- 	branch_block_stmt_2042/xx_xcritedgex_xix_xi_iq_err_calcx_xexit_PhiReq/phi_stmt_3568/phi_stmt_3568_sources/type_cast_3571/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_2042/xx_xcritedgex_xix_xi_iq_err_calcx_xexit_PhiReq/phi_stmt_3568/phi_stmt_3568_sources/type_cast_3571/SplitProtocol/Sample/ra
      -- 
    ra_19352_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3571_inst_ack_0, ack => cp_elements(2295)); -- 
    -- CP-element group 2296 transition  output  bypass 
    -- predecessors 989 
    -- successors 2297 
    -- members (2) 
      -- 	branch_block_stmt_2042/xx_xcritedgex_xix_xi_iq_err_calcx_xexit_PhiReq/phi_stmt_3568/phi_stmt_3568_sources/type_cast_3571/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_2042/xx_xcritedgex_xix_xi_iq_err_calcx_xexit_PhiReq/phi_stmt_3568/phi_stmt_3568_sources/type_cast_3571/SplitProtocol/Update/cr
      -- 
    cp_elements(2296) <= cp_elements(989);
    cr_19356_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2296), ack => type_cast_3571_inst_req_1); -- 
    -- CP-element group 2297 transition  input  bypass 
    -- predecessors 2296 
    -- successors 2298 
    -- members (2) 
      -- 	branch_block_stmt_2042/xx_xcritedgex_xix_xi_iq_err_calcx_xexit_PhiReq/phi_stmt_3568/phi_stmt_3568_sources/type_cast_3571/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_2042/xx_xcritedgex_xix_xi_iq_err_calcx_xexit_PhiReq/phi_stmt_3568/phi_stmt_3568_sources/type_cast_3571/SplitProtocol/Update/ca
      -- 
    ca_19357_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3571_inst_ack_1, ack => cp_elements(2297)); -- 
    -- CP-element group 2298 join  transition  output  bypass 
    -- predecessors 2295 2297 
    -- successors 2299 
    -- members (6) 
      -- 	branch_block_stmt_2042/xx_xcritedgex_xix_xi_iq_err_calcx_xexit_PhiReq/$exit
      -- 	branch_block_stmt_2042/xx_xcritedgex_xix_xi_iq_err_calcx_xexit_PhiReq/phi_stmt_3568/$exit
      -- 	branch_block_stmt_2042/xx_xcritedgex_xix_xi_iq_err_calcx_xexit_PhiReq/phi_stmt_3568/phi_stmt_3568_sources/$exit
      -- 	branch_block_stmt_2042/xx_xcritedgex_xix_xi_iq_err_calcx_xexit_PhiReq/phi_stmt_3568/phi_stmt_3568_sources/type_cast_3571/$exit
      -- 	branch_block_stmt_2042/xx_xcritedgex_xix_xi_iq_err_calcx_xexit_PhiReq/phi_stmt_3568/phi_stmt_3568_sources/type_cast_3571/SplitProtocol/$exit
      -- 	branch_block_stmt_2042/xx_xcritedgex_xix_xi_iq_err_calcx_xexit_PhiReq/phi_stmt_3568/phi_stmt_3568_req
      -- 
    cp_element_group_2298: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_2298"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(2295) & cp_elements(2297);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(2298), clk => clk, reset => reset); --
    end block;
    phi_stmt_3568_req_19358_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2298), ack => phi_stmt_3568_req_0); -- 
    -- CP-element group 2299 merge  place  bypass 
    -- predecessors 2293 2298 
    -- successors 2300 
    -- members (1) 
      -- 	branch_block_stmt_2042/merge_stmt_3567_PhiReqMerge
      -- 
    cp_elements(2299) <= OrReduce(cp_elements(2293) & cp_elements(2298));
    -- CP-element group 2300 transition  bypass 
    -- predecessors 2299 
    -- successors 2301 
    -- members (1) 
      -- 	branch_block_stmt_2042/merge_stmt_3567_PhiAck/$entry
      -- 
    cp_elements(2300) <= cp_elements(2299);
    -- CP-element group 2301 transition  place  input  bypass 
    -- predecessors 2300 
    -- successors 990 
    -- members (4) 
      -- 	branch_block_stmt_2042/assign_stmt_3580_to_assign_stmt_3603__entry__
      -- 	branch_block_stmt_2042/merge_stmt_3567__exit__
      -- 	branch_block_stmt_2042/merge_stmt_3567_PhiAck/$exit
      -- 	branch_block_stmt_2042/merge_stmt_3567_PhiAck/phi_stmt_3568_ack
      -- 
    phi_stmt_3568_ack_19363_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_3568_ack_0, ack => cp_elements(2301)); -- 
    -- CP-element group 2302 transition  bypass 
    -- predecessors 1027 
    -- successors 2304 
    -- members (4) 
      -- 	branch_block_stmt_2042/bb_56_bb_58_PhiReq/phi_stmt_3626/phi_stmt_3626_sources/type_cast_3629/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_2042/bb_56_bb_58_PhiReq/phi_stmt_3626/phi_stmt_3626_sources/type_cast_3629/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_2042/bb_56_bb_58_PhiReq/phi_stmt_3626/phi_stmt_3626_sources/type_cast_3629/SplitProtocol/Sample/rr
      -- 	branch_block_stmt_2042/bb_56_bb_58_PhiReq/phi_stmt_3626/phi_stmt_3626_sources/type_cast_3629/SplitProtocol/Sample/ra
      -- 
    cp_elements(2302) <= cp_elements(1027);
    -- CP-element group 2303 transition  bypass 
    -- predecessors 1027 
    -- successors 2304 
    -- members (4) 
      -- 	branch_block_stmt_2042/bb_56_bb_58_PhiReq/phi_stmt_3626/phi_stmt_3626_sources/type_cast_3629/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_2042/bb_56_bb_58_PhiReq/phi_stmt_3626/phi_stmt_3626_sources/type_cast_3629/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_2042/bb_56_bb_58_PhiReq/phi_stmt_3626/phi_stmt_3626_sources/type_cast_3629/SplitProtocol/Update/cr
      -- 	branch_block_stmt_2042/bb_56_bb_58_PhiReq/phi_stmt_3626/phi_stmt_3626_sources/type_cast_3629/SplitProtocol/Update/ca
      -- 
    cp_elements(2303) <= cp_elements(1027);
    -- CP-element group 2304 join  transition  output  bypass 
    -- predecessors 2302 2303 
    -- successors 2313 
    -- members (6) 
      -- 	branch_block_stmt_2042/bb_56_bb_58_PhiReq/$exit
      -- 	branch_block_stmt_2042/bb_56_bb_58_PhiReq/phi_stmt_3626/$exit
      -- 	branch_block_stmt_2042/bb_56_bb_58_PhiReq/phi_stmt_3626/phi_stmt_3626_sources/$exit
      -- 	branch_block_stmt_2042/bb_56_bb_58_PhiReq/phi_stmt_3626/phi_stmt_3626_sources/type_cast_3629/$exit
      -- 	branch_block_stmt_2042/bb_56_bb_58_PhiReq/phi_stmt_3626/phi_stmt_3626_sources/type_cast_3629/SplitProtocol/$exit
      -- 	branch_block_stmt_2042/bb_56_bb_58_PhiReq/phi_stmt_3626/phi_stmt_3626_req
      -- 
    cp_element_group_2304: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_2304"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(2302) & cp_elements(2303);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(2304), clk => clk, reset => reset); --
    end block;
    phi_stmt_3626_req_19413_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2304), ack => phi_stmt_3626_req_2); -- 
    -- CP-element group 2305 transition  output  bypass 
    -- predecessors 61 
    -- successors 2306 
    -- members (2) 
      -- 	branch_block_stmt_2042/bb_57_bb_58_PhiReq/phi_stmt_3626/phi_stmt_3626_sources/type_cast_3629/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_2042/bb_57_bb_58_PhiReq/phi_stmt_3626/phi_stmt_3626_sources/type_cast_3629/SplitProtocol/Sample/rr
      -- 
    cp_elements(2305) <= cp_elements(61);
    rr_19432_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2305), ack => type_cast_3629_inst_req_0); -- 
    -- CP-element group 2306 transition  input  bypass 
    -- predecessors 2305 
    -- successors 2309 
    -- members (2) 
      -- 	branch_block_stmt_2042/bb_57_bb_58_PhiReq/phi_stmt_3626/phi_stmt_3626_sources/type_cast_3629/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_2042/bb_57_bb_58_PhiReq/phi_stmt_3626/phi_stmt_3626_sources/type_cast_3629/SplitProtocol/Sample/ra
      -- 
    ra_19433_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3629_inst_ack_0, ack => cp_elements(2306)); -- 
    -- CP-element group 2307 transition  output  bypass 
    -- predecessors 61 
    -- successors 2308 
    -- members (2) 
      -- 	branch_block_stmt_2042/bb_57_bb_58_PhiReq/phi_stmt_3626/phi_stmt_3626_sources/type_cast_3629/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_2042/bb_57_bb_58_PhiReq/phi_stmt_3626/phi_stmt_3626_sources/type_cast_3629/SplitProtocol/Update/cr
      -- 
    cp_elements(2307) <= cp_elements(61);
    cr_19437_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2307), ack => type_cast_3629_inst_req_1); -- 
    -- CP-element group 2308 transition  input  bypass 
    -- predecessors 2307 
    -- successors 2309 
    -- members (2) 
      -- 	branch_block_stmt_2042/bb_57_bb_58_PhiReq/phi_stmt_3626/phi_stmt_3626_sources/type_cast_3629/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_2042/bb_57_bb_58_PhiReq/phi_stmt_3626/phi_stmt_3626_sources/type_cast_3629/SplitProtocol/Update/ca
      -- 
    ca_19438_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3629_inst_ack_1, ack => cp_elements(2308)); -- 
    -- CP-element group 2309 join  transition  output  bypass 
    -- predecessors 2306 2308 
    -- successors 2313 
    -- members (6) 
      -- 	branch_block_stmt_2042/bb_57_bb_58_PhiReq/$exit
      -- 	branch_block_stmt_2042/bb_57_bb_58_PhiReq/phi_stmt_3626/$exit
      -- 	branch_block_stmt_2042/bb_57_bb_58_PhiReq/phi_stmt_3626/phi_stmt_3626_sources/$exit
      -- 	branch_block_stmt_2042/bb_57_bb_58_PhiReq/phi_stmt_3626/phi_stmt_3626_sources/type_cast_3629/$exit
      -- 	branch_block_stmt_2042/bb_57_bb_58_PhiReq/phi_stmt_3626/phi_stmt_3626_sources/type_cast_3629/SplitProtocol/$exit
      -- 	branch_block_stmt_2042/bb_57_bb_58_PhiReq/phi_stmt_3626/phi_stmt_3626_req
      -- 
    cp_element_group_2309: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_2309"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(2306) & cp_elements(2308);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(2309), clk => clk, reset => reset); --
    end block;
    phi_stmt_3626_req_19439_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2309), ack => phi_stmt_3626_req_0); -- 
    -- CP-element group 2310 transition  bypass 
    -- predecessors 1015 
    -- successors 2312 
    -- members (4) 
      -- 	branch_block_stmt_2042/iq_err_calcx_xexit_bb_58_PhiReq/phi_stmt_3626/phi_stmt_3626_sources/type_cast_3629/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_2042/iq_err_calcx_xexit_bb_58_PhiReq/phi_stmt_3626/phi_stmt_3626_sources/type_cast_3629/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_2042/iq_err_calcx_xexit_bb_58_PhiReq/phi_stmt_3626/phi_stmt_3626_sources/type_cast_3629/SplitProtocol/Sample/rr
      -- 	branch_block_stmt_2042/iq_err_calcx_xexit_bb_58_PhiReq/phi_stmt_3626/phi_stmt_3626_sources/type_cast_3629/SplitProtocol/Sample/ra
      -- 
    cp_elements(2310) <= cp_elements(1015);
    -- CP-element group 2311 transition  bypass 
    -- predecessors 1015 
    -- successors 2312 
    -- members (4) 
      -- 	branch_block_stmt_2042/iq_err_calcx_xexit_bb_58_PhiReq/phi_stmt_3626/phi_stmt_3626_sources/type_cast_3629/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_2042/iq_err_calcx_xexit_bb_58_PhiReq/phi_stmt_3626/phi_stmt_3626_sources/type_cast_3629/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_2042/iq_err_calcx_xexit_bb_58_PhiReq/phi_stmt_3626/phi_stmt_3626_sources/type_cast_3629/SplitProtocol/Update/cr
      -- 	branch_block_stmt_2042/iq_err_calcx_xexit_bb_58_PhiReq/phi_stmt_3626/phi_stmt_3626_sources/type_cast_3629/SplitProtocol/Update/ca
      -- 
    cp_elements(2311) <= cp_elements(1015);
    -- CP-element group 2312 join  transition  output  bypass 
    -- predecessors 2310 2311 
    -- successors 2313 
    -- members (6) 
      -- 	branch_block_stmt_2042/iq_err_calcx_xexit_bb_58_PhiReq/$exit
      -- 	branch_block_stmt_2042/iq_err_calcx_xexit_bb_58_PhiReq/phi_stmt_3626/$exit
      -- 	branch_block_stmt_2042/iq_err_calcx_xexit_bb_58_PhiReq/phi_stmt_3626/phi_stmt_3626_sources/$exit
      -- 	branch_block_stmt_2042/iq_err_calcx_xexit_bb_58_PhiReq/phi_stmt_3626/phi_stmt_3626_sources/type_cast_3629/$exit
      -- 	branch_block_stmt_2042/iq_err_calcx_xexit_bb_58_PhiReq/phi_stmt_3626/phi_stmt_3626_sources/type_cast_3629/SplitProtocol/$exit
      -- 	branch_block_stmt_2042/iq_err_calcx_xexit_bb_58_PhiReq/phi_stmt_3626/phi_stmt_3626_req
      -- 
    cp_element_group_2312: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_2312"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(2310) & cp_elements(2311);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(2312), clk => clk, reset => reset); --
    end block;
    phi_stmt_3626_req_19465_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2312), ack => phi_stmt_3626_req_1); -- 
    -- CP-element group 2313 merge  place  bypass 
    -- predecessors 2304 2309 2312 
    -- successors 2314 
    -- members (1) 
      -- 	branch_block_stmt_2042/merge_stmt_3625_PhiReqMerge
      -- 
    cp_elements(2313) <= OrReduce(cp_elements(2304) & cp_elements(2309) & cp_elements(2312));
    -- CP-element group 2314 transition  bypass 
    -- predecessors 2313 
    -- successors 2315 
    -- members (1) 
      -- 	branch_block_stmt_2042/merge_stmt_3625_PhiAck/$entry
      -- 
    cp_elements(2314) <= cp_elements(2313);
    -- CP-element group 2315 transition  place  input  bypass 
    -- predecessors 2314 
    -- successors 1030 
    -- members (4) 
      -- 	branch_block_stmt_2042/assign_stmt_3642_to_assign_stmt_3653__entry__
      -- 	branch_block_stmt_2042/merge_stmt_3625__exit__
      -- 	branch_block_stmt_2042/merge_stmt_3625_PhiAck/$exit
      -- 	branch_block_stmt_2042/merge_stmt_3625_PhiAck/phi_stmt_3626_ack
      -- 
    phi_stmt_3626_ack_19470_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_3626_ack_0, ack => cp_elements(2315)); -- 
    -- CP-element group 2316 transition  bypass 
    -- predecessors 1047 
    -- successors 2318 
    -- members (4) 
      -- 	branch_block_stmt_2042/bb_58_xx_xthread_PhiReq/phi_stmt_3687/phi_stmt_3687_sources/type_cast_3690/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_2042/bb_58_xx_xthread_PhiReq/phi_stmt_3687/phi_stmt_3687_sources/type_cast_3690/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_2042/bb_58_xx_xthread_PhiReq/phi_stmt_3687/phi_stmt_3687_sources/type_cast_3690/SplitProtocol/Sample/rr
      -- 	branch_block_stmt_2042/bb_58_xx_xthread_PhiReq/phi_stmt_3687/phi_stmt_3687_sources/type_cast_3690/SplitProtocol/Sample/ra
      -- 
    cp_elements(2316) <= cp_elements(1047);
    -- CP-element group 2317 transition  bypass 
    -- predecessors 1047 
    -- successors 2318 
    -- members (4) 
      -- 	branch_block_stmt_2042/bb_58_xx_xthread_PhiReq/phi_stmt_3687/phi_stmt_3687_sources/type_cast_3690/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_2042/bb_58_xx_xthread_PhiReq/phi_stmt_3687/phi_stmt_3687_sources/type_cast_3690/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_2042/bb_58_xx_xthread_PhiReq/phi_stmt_3687/phi_stmt_3687_sources/type_cast_3690/SplitProtocol/Update/cr
      -- 	branch_block_stmt_2042/bb_58_xx_xthread_PhiReq/phi_stmt_3687/phi_stmt_3687_sources/type_cast_3690/SplitProtocol/Update/ca
      -- 
    cp_elements(2317) <= cp_elements(1047);
    -- CP-element group 2318 join  transition  output  bypass 
    -- predecessors 2316 2317 
    -- successors 2327 
    -- members (6) 
      -- 	branch_block_stmt_2042/bb_58_xx_xthread_PhiReq/$exit
      -- 	branch_block_stmt_2042/bb_58_xx_xthread_PhiReq/phi_stmt_3687/$exit
      -- 	branch_block_stmt_2042/bb_58_xx_xthread_PhiReq/phi_stmt_3687/phi_stmt_3687_sources/$exit
      -- 	branch_block_stmt_2042/bb_58_xx_xthread_PhiReq/phi_stmt_3687/phi_stmt_3687_sources/type_cast_3690/$exit
      -- 	branch_block_stmt_2042/bb_58_xx_xthread_PhiReq/phi_stmt_3687/phi_stmt_3687_sources/type_cast_3690/SplitProtocol/$exit
      -- 	branch_block_stmt_2042/bb_58_xx_xthread_PhiReq/phi_stmt_3687/phi_stmt_3687_req
      -- 
    cp_element_group_2318: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_2318"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(2316) & cp_elements(2317);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(2318), clk => clk, reset => reset); --
    end block;
    phi_stmt_3687_req_19524_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2318), ack => phi_stmt_3687_req_1); -- 
    -- CP-element group 2319 transition  bypass 
    -- predecessors 1059 
    -- successors 2321 
    -- members (4) 
      -- 	branch_block_stmt_2042/bb_59_xx_xthread_PhiReq/phi_stmt_3687/phi_stmt_3687_sources/type_cast_3690/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_2042/bb_59_xx_xthread_PhiReq/phi_stmt_3687/phi_stmt_3687_sources/type_cast_3690/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_2042/bb_59_xx_xthread_PhiReq/phi_stmt_3687/phi_stmt_3687_sources/type_cast_3690/SplitProtocol/Sample/rr
      -- 	branch_block_stmt_2042/bb_59_xx_xthread_PhiReq/phi_stmt_3687/phi_stmt_3687_sources/type_cast_3690/SplitProtocol/Sample/ra
      -- 
    cp_elements(2319) <= cp_elements(1059);
    -- CP-element group 2320 transition  bypass 
    -- predecessors 1059 
    -- successors 2321 
    -- members (4) 
      -- 	branch_block_stmt_2042/bb_59_xx_xthread_PhiReq/phi_stmt_3687/phi_stmt_3687_sources/type_cast_3690/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_2042/bb_59_xx_xthread_PhiReq/phi_stmt_3687/phi_stmt_3687_sources/type_cast_3690/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_2042/bb_59_xx_xthread_PhiReq/phi_stmt_3687/phi_stmt_3687_sources/type_cast_3690/SplitProtocol/Update/cr
      -- 	branch_block_stmt_2042/bb_59_xx_xthread_PhiReq/phi_stmt_3687/phi_stmt_3687_sources/type_cast_3690/SplitProtocol/Update/ca
      -- 
    cp_elements(2320) <= cp_elements(1059);
    -- CP-element group 2321 join  transition  output  bypass 
    -- predecessors 2319 2320 
    -- successors 2327 
    -- members (6) 
      -- 	branch_block_stmt_2042/bb_59_xx_xthread_PhiReq/$exit
      -- 	branch_block_stmt_2042/bb_59_xx_xthread_PhiReq/phi_stmt_3687/$exit
      -- 	branch_block_stmt_2042/bb_59_xx_xthread_PhiReq/phi_stmt_3687/phi_stmt_3687_sources/$exit
      -- 	branch_block_stmt_2042/bb_59_xx_xthread_PhiReq/phi_stmt_3687/phi_stmt_3687_sources/type_cast_3690/$exit
      -- 	branch_block_stmt_2042/bb_59_xx_xthread_PhiReq/phi_stmt_3687/phi_stmt_3687_sources/type_cast_3690/SplitProtocol/$exit
      -- 	branch_block_stmt_2042/bb_59_xx_xthread_PhiReq/phi_stmt_3687/phi_stmt_3687_req
      -- 
    cp_element_group_2321: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_2321"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(2319) & cp_elements(2320);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(2321), clk => clk, reset => reset); --
    end block;
    phi_stmt_3687_req_19550_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2321), ack => phi_stmt_3687_req_2); -- 
    -- CP-element group 2322 transition  output  bypass 
    -- predecessors 1073 
    -- successors 2323 
    -- members (2) 
      -- 	branch_block_stmt_2042/bb_60_xx_xthread_PhiReq/phi_stmt_3687/phi_stmt_3687_sources/type_cast_3690/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_2042/bb_60_xx_xthread_PhiReq/phi_stmt_3687/phi_stmt_3687_sources/type_cast_3690/SplitProtocol/Sample/rr
      -- 
    cp_elements(2322) <= cp_elements(1073);
    rr_19569_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2322), ack => type_cast_3690_inst_req_0); -- 
    -- CP-element group 2323 transition  input  bypass 
    -- predecessors 2322 
    -- successors 2326 
    -- members (2) 
      -- 	branch_block_stmt_2042/bb_60_xx_xthread_PhiReq/phi_stmt_3687/phi_stmt_3687_sources/type_cast_3690/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_2042/bb_60_xx_xthread_PhiReq/phi_stmt_3687/phi_stmt_3687_sources/type_cast_3690/SplitProtocol/Sample/ra
      -- 
    ra_19570_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3690_inst_ack_0, ack => cp_elements(2323)); -- 
    -- CP-element group 2324 transition  output  bypass 
    -- predecessors 1073 
    -- successors 2325 
    -- members (2) 
      -- 	branch_block_stmt_2042/bb_60_xx_xthread_PhiReq/phi_stmt_3687/phi_stmt_3687_sources/type_cast_3690/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_2042/bb_60_xx_xthread_PhiReq/phi_stmt_3687/phi_stmt_3687_sources/type_cast_3690/SplitProtocol/Update/cr
      -- 
    cp_elements(2324) <= cp_elements(1073);
    cr_19574_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2324), ack => type_cast_3690_inst_req_1); -- 
    -- CP-element group 2325 transition  input  bypass 
    -- predecessors 2324 
    -- successors 2326 
    -- members (2) 
      -- 	branch_block_stmt_2042/bb_60_xx_xthread_PhiReq/phi_stmt_3687/phi_stmt_3687_sources/type_cast_3690/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_2042/bb_60_xx_xthread_PhiReq/phi_stmt_3687/phi_stmt_3687_sources/type_cast_3690/SplitProtocol/Update/ca
      -- 
    ca_19575_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3690_inst_ack_1, ack => cp_elements(2325)); -- 
    -- CP-element group 2326 join  transition  output  bypass 
    -- predecessors 2323 2325 
    -- successors 2327 
    -- members (6) 
      -- 	branch_block_stmt_2042/bb_60_xx_xthread_PhiReq/$exit
      -- 	branch_block_stmt_2042/bb_60_xx_xthread_PhiReq/phi_stmt_3687/$exit
      -- 	branch_block_stmt_2042/bb_60_xx_xthread_PhiReq/phi_stmt_3687/phi_stmt_3687_sources/$exit
      -- 	branch_block_stmt_2042/bb_60_xx_xthread_PhiReq/phi_stmt_3687/phi_stmt_3687_sources/type_cast_3690/$exit
      -- 	branch_block_stmt_2042/bb_60_xx_xthread_PhiReq/phi_stmt_3687/phi_stmt_3687_sources/type_cast_3690/SplitProtocol/$exit
      -- 	branch_block_stmt_2042/bb_60_xx_xthread_PhiReq/phi_stmt_3687/phi_stmt_3687_req
      -- 
    cp_element_group_2326: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_2326"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(2323) & cp_elements(2325);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(2326), clk => clk, reset => reset); --
    end block;
    phi_stmt_3687_req_19576_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2326), ack => phi_stmt_3687_req_0); -- 
    -- CP-element group 2327 merge  place  bypass 
    -- predecessors 2318 2321 2326 
    -- successors 2328 
    -- members (1) 
      -- 	branch_block_stmt_2042/merge_stmt_3686_PhiReqMerge
      -- 
    cp_elements(2327) <= OrReduce(cp_elements(2318) & cp_elements(2321) & cp_elements(2326));
    -- CP-element group 2328 transition  bypass 
    -- predecessors 2327 
    -- successors 2329 
    -- members (1) 
      -- 	branch_block_stmt_2042/merge_stmt_3686_PhiAck/$entry
      -- 
    cp_elements(2328) <= cp_elements(2327);
    -- CP-element group 2329 transition  input  bypass 
    -- predecessors 2328 
    -- successors 64 
    -- members (2) 
      -- 	branch_block_stmt_2042/merge_stmt_3686_PhiAck/$exit
      -- 	branch_block_stmt_2042/merge_stmt_3686_PhiAck/phi_stmt_3687_ack
      -- 
    phi_stmt_3687_ack_19581_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_3687_ack_0, ack => cp_elements(2329)); -- 
    -- CP-element group 2330 fork  transition  bypass 
    -- predecessors 1148 
    -- successors 2331 2343 
    -- members (1) 
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xi_bbx_xnph7x_xix_xi_PhiReq/$entry
      -- 
    cp_elements(2330) <= cp_elements(1148);
    -- CP-element group 2331 fork  transition  bypass 
    -- predecessors 2330 
    -- successors 2332 2338 
    -- members (2) 
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xi_bbx_xnph7x_xix_xi_PhiReq/phi_stmt_3722/$entry
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xi_bbx_xnph7x_xix_xi_PhiReq/phi_stmt_3722/phi_stmt_3722_sources/$entry
      -- 
    cp_elements(2331) <= cp_elements(2330);
    -- CP-element group 2332 fork  transition  bypass 
    -- predecessors 2331 
    -- successors 2333 2335 
    -- members (2) 
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xi_bbx_xnph7x_xix_xi_PhiReq/phi_stmt_3722/phi_stmt_3722_sources/type_cast_3725/$entry
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xi_bbx_xnph7x_xix_xi_PhiReq/phi_stmt_3722/phi_stmt_3722_sources/type_cast_3725/SplitProtocol/$entry
      -- 
    cp_elements(2332) <= cp_elements(2331);
    -- CP-element group 2333 transition  output  bypass 
    -- predecessors 2332 
    -- successors 2334 
    -- members (2) 
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xi_bbx_xnph7x_xix_xi_PhiReq/phi_stmt_3722/phi_stmt_3722_sources/type_cast_3725/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xi_bbx_xnph7x_xix_xi_PhiReq/phi_stmt_3722/phi_stmt_3722_sources/type_cast_3725/SplitProtocol/Sample/rr
      -- 
    cp_elements(2333) <= cp_elements(2332);
    rr_19600_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2333), ack => type_cast_3725_inst_req_0); -- 
    -- CP-element group 2334 transition  input  bypass 
    -- predecessors 2333 
    -- successors 2337 
    -- members (2) 
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xi_bbx_xnph7x_xix_xi_PhiReq/phi_stmt_3722/phi_stmt_3722_sources/type_cast_3725/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xi_bbx_xnph7x_xix_xi_PhiReq/phi_stmt_3722/phi_stmt_3722_sources/type_cast_3725/SplitProtocol/Sample/ra
      -- 
    ra_19601_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3725_inst_ack_0, ack => cp_elements(2334)); -- 
    -- CP-element group 2335 transition  output  bypass 
    -- predecessors 2332 
    -- successors 2336 
    -- members (2) 
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xi_bbx_xnph7x_xix_xi_PhiReq/phi_stmt_3722/phi_stmt_3722_sources/type_cast_3725/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xi_bbx_xnph7x_xix_xi_PhiReq/phi_stmt_3722/phi_stmt_3722_sources/type_cast_3725/SplitProtocol/Update/cr
      -- 
    cp_elements(2335) <= cp_elements(2332);
    cr_19605_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2335), ack => type_cast_3725_inst_req_1); -- 
    -- CP-element group 2336 transition  input  bypass 
    -- predecessors 2335 
    -- successors 2337 
    -- members (2) 
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xi_bbx_xnph7x_xix_xi_PhiReq/phi_stmt_3722/phi_stmt_3722_sources/type_cast_3725/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xi_bbx_xnph7x_xix_xi_PhiReq/phi_stmt_3722/phi_stmt_3722_sources/type_cast_3725/SplitProtocol/Update/ca
      -- 
    ca_19606_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3725_inst_ack_1, ack => cp_elements(2336)); -- 
    -- CP-element group 2337 join  transition  bypass 
    -- predecessors 2334 2336 
    -- successors 2342 
    -- members (2) 
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xi_bbx_xnph7x_xix_xi_PhiReq/phi_stmt_3722/phi_stmt_3722_sources/type_cast_3725/$exit
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xi_bbx_xnph7x_xix_xi_PhiReq/phi_stmt_3722/phi_stmt_3722_sources/type_cast_3725/SplitProtocol/$exit
      -- 
    cp_element_group_2337: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_2337"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(2334) & cp_elements(2336);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(2337), clk => clk, reset => reset); --
    end block;
    -- CP-element group 2338 fork  transition  bypass 
    -- predecessors 2331 
    -- successors 2339 2340 
    -- members (2) 
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xi_bbx_xnph7x_xix_xi_PhiReq/phi_stmt_3722/phi_stmt_3722_sources/type_cast_3727/$entry
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xi_bbx_xnph7x_xix_xi_PhiReq/phi_stmt_3722/phi_stmt_3722_sources/type_cast_3727/SplitProtocol/$entry
      -- 
    cp_elements(2338) <= cp_elements(2331);
    -- CP-element group 2339 transition  bypass 
    -- predecessors 2338 
    -- successors 2341 
    -- members (4) 
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xi_bbx_xnph7x_xix_xi_PhiReq/phi_stmt_3722/phi_stmt_3722_sources/type_cast_3727/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xi_bbx_xnph7x_xix_xi_PhiReq/phi_stmt_3722/phi_stmt_3722_sources/type_cast_3727/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xi_bbx_xnph7x_xix_xi_PhiReq/phi_stmt_3722/phi_stmt_3722_sources/type_cast_3727/SplitProtocol/Sample/rr
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xi_bbx_xnph7x_xix_xi_PhiReq/phi_stmt_3722/phi_stmt_3722_sources/type_cast_3727/SplitProtocol/Sample/ra
      -- 
    cp_elements(2339) <= cp_elements(2338);
    -- CP-element group 2340 transition  bypass 
    -- predecessors 2338 
    -- successors 2341 
    -- members (4) 
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xi_bbx_xnph7x_xix_xi_PhiReq/phi_stmt_3722/phi_stmt_3722_sources/type_cast_3727/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xi_bbx_xnph7x_xix_xi_PhiReq/phi_stmt_3722/phi_stmt_3722_sources/type_cast_3727/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xi_bbx_xnph7x_xix_xi_PhiReq/phi_stmt_3722/phi_stmt_3722_sources/type_cast_3727/SplitProtocol/Update/cr
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xi_bbx_xnph7x_xix_xi_PhiReq/phi_stmt_3722/phi_stmt_3722_sources/type_cast_3727/SplitProtocol/Update/ca
      -- 
    cp_elements(2340) <= cp_elements(2338);
    -- CP-element group 2341 join  transition  bypass 
    -- predecessors 2339 2340 
    -- successors 2342 
    -- members (2) 
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xi_bbx_xnph7x_xix_xi_PhiReq/phi_stmt_3722/phi_stmt_3722_sources/type_cast_3727/$exit
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xi_bbx_xnph7x_xix_xi_PhiReq/phi_stmt_3722/phi_stmt_3722_sources/type_cast_3727/SplitProtocol/$exit
      -- 
    cp_element_group_2341: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_2341"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(2339) & cp_elements(2340);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(2341), clk => clk, reset => reset); --
    end block;
    -- CP-element group 2342 join  transition  output  bypass 
    -- predecessors 2337 2341 
    -- successors 2349 
    -- members (3) 
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xi_bbx_xnph7x_xix_xi_PhiReq/phi_stmt_3722/$exit
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xi_bbx_xnph7x_xix_xi_PhiReq/phi_stmt_3722/phi_stmt_3722_sources/$exit
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xi_bbx_xnph7x_xix_xi_PhiReq/phi_stmt_3722/phi_stmt_3722_req
      -- 
    cp_element_group_2342: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_2342"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(2337) & cp_elements(2341);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(2342), clk => clk, reset => reset); --
    end block;
    phi_stmt_3722_req_19623_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2342), ack => phi_stmt_3722_req_0); -- 
    -- CP-element group 2343 fork  transition  bypass 
    -- predecessors 2330 
    -- successors 2344 2346 
    -- members (4) 
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xi_bbx_xnph7x_xix_xi_PhiReq/phi_stmt_3728/$entry
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xi_bbx_xnph7x_xix_xi_PhiReq/phi_stmt_3728/phi_stmt_3728_sources/$entry
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xi_bbx_xnph7x_xix_xi_PhiReq/phi_stmt_3728/phi_stmt_3728_sources/type_cast_3731/$entry
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xi_bbx_xnph7x_xix_xi_PhiReq/phi_stmt_3728/phi_stmt_3728_sources/type_cast_3731/SplitProtocol/$entry
      -- 
    cp_elements(2343) <= cp_elements(2330);
    -- CP-element group 2344 transition  output  bypass 
    -- predecessors 2343 
    -- successors 2345 
    -- members (2) 
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xi_bbx_xnph7x_xix_xi_PhiReq/phi_stmt_3728/phi_stmt_3728_sources/type_cast_3731/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xi_bbx_xnph7x_xix_xi_PhiReq/phi_stmt_3728/phi_stmt_3728_sources/type_cast_3731/SplitProtocol/Sample/rr
      -- 
    cp_elements(2344) <= cp_elements(2343);
    rr_19639_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2344), ack => type_cast_3731_inst_req_0); -- 
    -- CP-element group 2345 transition  input  bypass 
    -- predecessors 2344 
    -- successors 2348 
    -- members (2) 
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xi_bbx_xnph7x_xix_xi_PhiReq/phi_stmt_3728/phi_stmt_3728_sources/type_cast_3731/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xi_bbx_xnph7x_xix_xi_PhiReq/phi_stmt_3728/phi_stmt_3728_sources/type_cast_3731/SplitProtocol/Sample/ra
      -- 
    ra_19640_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3731_inst_ack_0, ack => cp_elements(2345)); -- 
    -- CP-element group 2346 transition  output  bypass 
    -- predecessors 2343 
    -- successors 2347 
    -- members (2) 
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xi_bbx_xnph7x_xix_xi_PhiReq/phi_stmt_3728/phi_stmt_3728_sources/type_cast_3731/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xi_bbx_xnph7x_xix_xi_PhiReq/phi_stmt_3728/phi_stmt_3728_sources/type_cast_3731/SplitProtocol/Update/cr
      -- 
    cp_elements(2346) <= cp_elements(2343);
    cr_19644_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2346), ack => type_cast_3731_inst_req_1); -- 
    -- CP-element group 2347 transition  input  bypass 
    -- predecessors 2346 
    -- successors 2348 
    -- members (2) 
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xi_bbx_xnph7x_xix_xi_PhiReq/phi_stmt_3728/phi_stmt_3728_sources/type_cast_3731/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xi_bbx_xnph7x_xix_xi_PhiReq/phi_stmt_3728/phi_stmt_3728_sources/type_cast_3731/SplitProtocol/Update/ca
      -- 
    ca_19645_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3731_inst_ack_1, ack => cp_elements(2347)); -- 
    -- CP-element group 2348 join  transition  output  bypass 
    -- predecessors 2345 2347 
    -- successors 2349 
    -- members (5) 
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xi_bbx_xnph7x_xix_xi_PhiReq/phi_stmt_3728/$exit
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xi_bbx_xnph7x_xix_xi_PhiReq/phi_stmt_3728/phi_stmt_3728_sources/$exit
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xi_bbx_xnph7x_xix_xi_PhiReq/phi_stmt_3728/phi_stmt_3728_sources/type_cast_3731/$exit
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xi_bbx_xnph7x_xix_xi_PhiReq/phi_stmt_3728/phi_stmt_3728_sources/type_cast_3731/SplitProtocol/$exit
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xi_bbx_xnph7x_xix_xi_PhiReq/phi_stmt_3728/phi_stmt_3728_req
      -- 
    cp_element_group_2348: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_2348"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(2345) & cp_elements(2347);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(2348), clk => clk, reset => reset); --
    end block;
    phi_stmt_3728_req_19646_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2348), ack => phi_stmt_3728_req_0); -- 
    -- CP-element group 2349 join  transition  bypass 
    -- predecessors 2342 2348 
    -- successors 2368 
    -- members (1) 
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xi_bbx_xnph7x_xix_xi_PhiReq/$exit
      -- 
    cp_element_group_2349: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_2349"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(2342) & cp_elements(2348);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(2349), clk => clk, reset => reset); --
    end block;
    -- CP-element group 2350 fork  transition  bypass 
    -- predecessors 1087 
    -- successors 2351 2363 
    -- members (1) 
      -- 	branch_block_stmt_2042/xx_xthread_bbx_xnph7x_xix_xi_PhiReq/$entry
      -- 
    cp_elements(2350) <= cp_elements(1087);
    -- CP-element group 2351 fork  transition  bypass 
    -- predecessors 2350 
    -- successors 2352 2356 
    -- members (2) 
      -- 	branch_block_stmt_2042/xx_xthread_bbx_xnph7x_xix_xi_PhiReq/phi_stmt_3722/$entry
      -- 	branch_block_stmt_2042/xx_xthread_bbx_xnph7x_xix_xi_PhiReq/phi_stmt_3722/phi_stmt_3722_sources/$entry
      -- 
    cp_elements(2351) <= cp_elements(2350);
    -- CP-element group 2352 fork  transition  bypass 
    -- predecessors 2351 
    -- successors 2353 2354 
    -- members (2) 
      -- 	branch_block_stmt_2042/xx_xthread_bbx_xnph7x_xix_xi_PhiReq/phi_stmt_3722/phi_stmt_3722_sources/type_cast_3725/$entry
      -- 	branch_block_stmt_2042/xx_xthread_bbx_xnph7x_xix_xi_PhiReq/phi_stmt_3722/phi_stmt_3722_sources/type_cast_3725/SplitProtocol/$entry
      -- 
    cp_elements(2352) <= cp_elements(2351);
    -- CP-element group 2353 transition  bypass 
    -- predecessors 2352 
    -- successors 2355 
    -- members (4) 
      -- 	branch_block_stmt_2042/xx_xthread_bbx_xnph7x_xix_xi_PhiReq/phi_stmt_3722/phi_stmt_3722_sources/type_cast_3725/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_2042/xx_xthread_bbx_xnph7x_xix_xi_PhiReq/phi_stmt_3722/phi_stmt_3722_sources/type_cast_3725/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_2042/xx_xthread_bbx_xnph7x_xix_xi_PhiReq/phi_stmt_3722/phi_stmt_3722_sources/type_cast_3725/SplitProtocol/Sample/rr
      -- 	branch_block_stmt_2042/xx_xthread_bbx_xnph7x_xix_xi_PhiReq/phi_stmt_3722/phi_stmt_3722_sources/type_cast_3725/SplitProtocol/Sample/ra
      -- 
    cp_elements(2353) <= cp_elements(2352);
    -- CP-element group 2354 transition  bypass 
    -- predecessors 2352 
    -- successors 2355 
    -- members (4) 
      -- 	branch_block_stmt_2042/xx_xthread_bbx_xnph7x_xix_xi_PhiReq/phi_stmt_3722/phi_stmt_3722_sources/type_cast_3725/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_2042/xx_xthread_bbx_xnph7x_xix_xi_PhiReq/phi_stmt_3722/phi_stmt_3722_sources/type_cast_3725/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_2042/xx_xthread_bbx_xnph7x_xix_xi_PhiReq/phi_stmt_3722/phi_stmt_3722_sources/type_cast_3725/SplitProtocol/Update/cr
      -- 	branch_block_stmt_2042/xx_xthread_bbx_xnph7x_xix_xi_PhiReq/phi_stmt_3722/phi_stmt_3722_sources/type_cast_3725/SplitProtocol/Update/ca
      -- 
    cp_elements(2354) <= cp_elements(2352);
    -- CP-element group 2355 join  transition  bypass 
    -- predecessors 2353 2354 
    -- successors 2362 
    -- members (2) 
      -- 	branch_block_stmt_2042/xx_xthread_bbx_xnph7x_xix_xi_PhiReq/phi_stmt_3722/phi_stmt_3722_sources/type_cast_3725/$exit
      -- 	branch_block_stmt_2042/xx_xthread_bbx_xnph7x_xix_xi_PhiReq/phi_stmt_3722/phi_stmt_3722_sources/type_cast_3725/SplitProtocol/$exit
      -- 
    cp_element_group_2355: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_2355"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(2353) & cp_elements(2354);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(2355), clk => clk, reset => reset); --
    end block;
    -- CP-element group 2356 fork  transition  bypass 
    -- predecessors 2351 
    -- successors 2357 2359 
    -- members (2) 
      -- 	branch_block_stmt_2042/xx_xthread_bbx_xnph7x_xix_xi_PhiReq/phi_stmt_3722/phi_stmt_3722_sources/type_cast_3727/$entry
      -- 	branch_block_stmt_2042/xx_xthread_bbx_xnph7x_xix_xi_PhiReq/phi_stmt_3722/phi_stmt_3722_sources/type_cast_3727/SplitProtocol/$entry
      -- 
    cp_elements(2356) <= cp_elements(2351);
    -- CP-element group 2357 transition  output  bypass 
    -- predecessors 2356 
    -- successors 2358 
    -- members (2) 
      -- 	branch_block_stmt_2042/xx_xthread_bbx_xnph7x_xix_xi_PhiReq/phi_stmt_3722/phi_stmt_3722_sources/type_cast_3727/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_2042/xx_xthread_bbx_xnph7x_xix_xi_PhiReq/phi_stmt_3722/phi_stmt_3722_sources/type_cast_3727/SplitProtocol/Sample/rr
      -- 
    cp_elements(2357) <= cp_elements(2356);
    rr_19681_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2357), ack => type_cast_3727_inst_req_0); -- 
    -- CP-element group 2358 transition  input  bypass 
    -- predecessors 2357 
    -- successors 2361 
    -- members (2) 
      -- 	branch_block_stmt_2042/xx_xthread_bbx_xnph7x_xix_xi_PhiReq/phi_stmt_3722/phi_stmt_3722_sources/type_cast_3727/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_2042/xx_xthread_bbx_xnph7x_xix_xi_PhiReq/phi_stmt_3722/phi_stmt_3722_sources/type_cast_3727/SplitProtocol/Sample/ra
      -- 
    ra_19682_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3727_inst_ack_0, ack => cp_elements(2358)); -- 
    -- CP-element group 2359 transition  output  bypass 
    -- predecessors 2356 
    -- successors 2360 
    -- members (2) 
      -- 	branch_block_stmt_2042/xx_xthread_bbx_xnph7x_xix_xi_PhiReq/phi_stmt_3722/phi_stmt_3722_sources/type_cast_3727/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_2042/xx_xthread_bbx_xnph7x_xix_xi_PhiReq/phi_stmt_3722/phi_stmt_3722_sources/type_cast_3727/SplitProtocol/Update/cr
      -- 
    cp_elements(2359) <= cp_elements(2356);
    cr_19686_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2359), ack => type_cast_3727_inst_req_1); -- 
    -- CP-element group 2360 transition  input  bypass 
    -- predecessors 2359 
    -- successors 2361 
    -- members (2) 
      -- 	branch_block_stmt_2042/xx_xthread_bbx_xnph7x_xix_xi_PhiReq/phi_stmt_3722/phi_stmt_3722_sources/type_cast_3727/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_2042/xx_xthread_bbx_xnph7x_xix_xi_PhiReq/phi_stmt_3722/phi_stmt_3722_sources/type_cast_3727/SplitProtocol/Update/ca
      -- 
    ca_19687_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3727_inst_ack_1, ack => cp_elements(2360)); -- 
    -- CP-element group 2361 join  transition  bypass 
    -- predecessors 2358 2360 
    -- successors 2362 
    -- members (2) 
      -- 	branch_block_stmt_2042/xx_xthread_bbx_xnph7x_xix_xi_PhiReq/phi_stmt_3722/phi_stmt_3722_sources/type_cast_3727/$exit
      -- 	branch_block_stmt_2042/xx_xthread_bbx_xnph7x_xix_xi_PhiReq/phi_stmt_3722/phi_stmt_3722_sources/type_cast_3727/SplitProtocol/$exit
      -- 
    cp_element_group_2361: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_2361"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(2358) & cp_elements(2360);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(2361), clk => clk, reset => reset); --
    end block;
    -- CP-element group 2362 join  transition  output  bypass 
    -- predecessors 2355 2361 
    -- successors 2367 
    -- members (3) 
      -- 	branch_block_stmt_2042/xx_xthread_bbx_xnph7x_xix_xi_PhiReq/phi_stmt_3722/$exit
      -- 	branch_block_stmt_2042/xx_xthread_bbx_xnph7x_xix_xi_PhiReq/phi_stmt_3722/phi_stmt_3722_sources/$exit
      -- 	branch_block_stmt_2042/xx_xthread_bbx_xnph7x_xix_xi_PhiReq/phi_stmt_3722/phi_stmt_3722_req
      -- 
    cp_element_group_2362: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_2362"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(2355) & cp_elements(2361);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(2362), clk => clk, reset => reset); --
    end block;
    phi_stmt_3722_req_19688_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2362), ack => phi_stmt_3722_req_1); -- 
    -- CP-element group 2363 fork  transition  bypass 
    -- predecessors 2350 
    -- successors 2364 2365 
    -- members (4) 
      -- 	branch_block_stmt_2042/xx_xthread_bbx_xnph7x_xix_xi_PhiReq/phi_stmt_3728/$entry
      -- 	branch_block_stmt_2042/xx_xthread_bbx_xnph7x_xix_xi_PhiReq/phi_stmt_3728/phi_stmt_3728_sources/$entry
      -- 	branch_block_stmt_2042/xx_xthread_bbx_xnph7x_xix_xi_PhiReq/phi_stmt_3728/phi_stmt_3728_sources/type_cast_3731/$entry
      -- 	branch_block_stmt_2042/xx_xthread_bbx_xnph7x_xix_xi_PhiReq/phi_stmt_3728/phi_stmt_3728_sources/type_cast_3731/SplitProtocol/$entry
      -- 
    cp_elements(2363) <= cp_elements(2350);
    -- CP-element group 2364 transition  bypass 
    -- predecessors 2363 
    -- successors 2366 
    -- members (4) 
      -- 	branch_block_stmt_2042/xx_xthread_bbx_xnph7x_xix_xi_PhiReq/phi_stmt_3728/phi_stmt_3728_sources/type_cast_3731/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_2042/xx_xthread_bbx_xnph7x_xix_xi_PhiReq/phi_stmt_3728/phi_stmt_3728_sources/type_cast_3731/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_2042/xx_xthread_bbx_xnph7x_xix_xi_PhiReq/phi_stmt_3728/phi_stmt_3728_sources/type_cast_3731/SplitProtocol/Sample/rr
      -- 	branch_block_stmt_2042/xx_xthread_bbx_xnph7x_xix_xi_PhiReq/phi_stmt_3728/phi_stmt_3728_sources/type_cast_3731/SplitProtocol/Sample/ra
      -- 
    cp_elements(2364) <= cp_elements(2363);
    -- CP-element group 2365 transition  bypass 
    -- predecessors 2363 
    -- successors 2366 
    -- members (4) 
      -- 	branch_block_stmt_2042/xx_xthread_bbx_xnph7x_xix_xi_PhiReq/phi_stmt_3728/phi_stmt_3728_sources/type_cast_3731/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_2042/xx_xthread_bbx_xnph7x_xix_xi_PhiReq/phi_stmt_3728/phi_stmt_3728_sources/type_cast_3731/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_2042/xx_xthread_bbx_xnph7x_xix_xi_PhiReq/phi_stmt_3728/phi_stmt_3728_sources/type_cast_3731/SplitProtocol/Update/cr
      -- 	branch_block_stmt_2042/xx_xthread_bbx_xnph7x_xix_xi_PhiReq/phi_stmt_3728/phi_stmt_3728_sources/type_cast_3731/SplitProtocol/Update/ca
      -- 
    cp_elements(2365) <= cp_elements(2363);
    -- CP-element group 2366 join  transition  output  bypass 
    -- predecessors 2364 2365 
    -- successors 2367 
    -- members (5) 
      -- 	branch_block_stmt_2042/xx_xthread_bbx_xnph7x_xix_xi_PhiReq/phi_stmt_3728/$exit
      -- 	branch_block_stmt_2042/xx_xthread_bbx_xnph7x_xix_xi_PhiReq/phi_stmt_3728/phi_stmt_3728_sources/$exit
      -- 	branch_block_stmt_2042/xx_xthread_bbx_xnph7x_xix_xi_PhiReq/phi_stmt_3728/phi_stmt_3728_sources/type_cast_3731/$exit
      -- 	branch_block_stmt_2042/xx_xthread_bbx_xnph7x_xix_xi_PhiReq/phi_stmt_3728/phi_stmt_3728_sources/type_cast_3731/SplitProtocol/$exit
      -- 	branch_block_stmt_2042/xx_xthread_bbx_xnph7x_xix_xi_PhiReq/phi_stmt_3728/phi_stmt_3728_req
      -- 
    cp_element_group_2366: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_2366"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(2364) & cp_elements(2365);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(2366), clk => clk, reset => reset); --
    end block;
    phi_stmt_3728_req_19711_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2366), ack => phi_stmt_3728_req_1); -- 
    -- CP-element group 2367 join  transition  bypass 
    -- predecessors 2362 2366 
    -- successors 2368 
    -- members (1) 
      -- 	branch_block_stmt_2042/xx_xthread_bbx_xnph7x_xix_xi_PhiReq/$exit
      -- 
    cp_element_group_2367: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_2367"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(2362) & cp_elements(2366);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(2367), clk => clk, reset => reset); --
    end block;
    -- CP-element group 2368 merge  place  bypass 
    -- predecessors 2349 2367 
    -- successors 2369 
    -- members (1) 
      -- 	branch_block_stmt_2042/merge_stmt_3721_PhiReqMerge
      -- 
    cp_elements(2368) <= OrReduce(cp_elements(2349) & cp_elements(2367));
    -- CP-element group 2369 fork  transition  bypass 
    -- predecessors 2368 
    -- successors 2370 2371 
    -- members (1) 
      -- 	branch_block_stmt_2042/merge_stmt_3721_PhiAck/$entry
      -- 
    cp_elements(2369) <= cp_elements(2368);
    -- CP-element group 2370 transition  input  bypass 
    -- predecessors 2369 
    -- successors 2372 
    -- members (1) 
      -- 	branch_block_stmt_2042/merge_stmt_3721_PhiAck/phi_stmt_3722_ack
      -- 
    phi_stmt_3722_ack_19716_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_3722_ack_0, ack => cp_elements(2370)); -- 
    -- CP-element group 2371 transition  input  bypass 
    -- predecessors 2369 
    -- successors 2372 
    -- members (1) 
      -- 	branch_block_stmt_2042/merge_stmt_3721_PhiAck/phi_stmt_3728_ack
      -- 
    phi_stmt_3728_ack_19717_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_3728_ack_0, ack => cp_elements(2371)); -- 
    -- CP-element group 2372 join  transition  bypass 
    -- predecessors 2370 2371 
    -- successors 65 
    -- members (1) 
      -- 	branch_block_stmt_2042/merge_stmt_3721_PhiAck/$exit
      -- 
    cp_element_group_2372: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_2372"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(2370) & cp_elements(2371);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(2372), clk => clk, reset => reset); --
    end block;
    -- CP-element group 2373 fork  transition  bypass 
    -- predecessors 1122 
    -- successors 2374 2380 
    -- members (1) 
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xi_bbx_xnphx_xix_xi_PhiReq/$entry
      -- 
    cp_elements(2373) <= cp_elements(1122);
    -- CP-element group 2374 fork  transition  bypass 
    -- predecessors 2373 
    -- successors 2375 2377 
    -- members (4) 
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xi_bbx_xnphx_xix_xi_PhiReq/phi_stmt_3757/$entry
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xi_bbx_xnphx_xix_xi_PhiReq/phi_stmt_3757/phi_stmt_3757_sources/$entry
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xi_bbx_xnphx_xix_xi_PhiReq/phi_stmt_3757/phi_stmt_3757_sources/type_cast_3760/$entry
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xi_bbx_xnphx_xix_xi_PhiReq/phi_stmt_3757/phi_stmt_3757_sources/type_cast_3760/SplitProtocol/$entry
      -- 
    cp_elements(2374) <= cp_elements(2373);
    -- CP-element group 2375 transition  output  bypass 
    -- predecessors 2374 
    -- successors 2376 
    -- members (2) 
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xi_bbx_xnphx_xix_xi_PhiReq/phi_stmt_3757/phi_stmt_3757_sources/type_cast_3760/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xi_bbx_xnphx_xix_xi_PhiReq/phi_stmt_3757/phi_stmt_3757_sources/type_cast_3760/SplitProtocol/Sample/rr
      -- 
    cp_elements(2375) <= cp_elements(2374);
    rr_19748_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2375), ack => type_cast_3760_inst_req_0); -- 
    -- CP-element group 2376 transition  input  bypass 
    -- predecessors 2375 
    -- successors 2379 
    -- members (2) 
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xi_bbx_xnphx_xix_xi_PhiReq/phi_stmt_3757/phi_stmt_3757_sources/type_cast_3760/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xi_bbx_xnphx_xix_xi_PhiReq/phi_stmt_3757/phi_stmt_3757_sources/type_cast_3760/SplitProtocol/Sample/ra
      -- 
    ra_19749_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3760_inst_ack_0, ack => cp_elements(2376)); -- 
    -- CP-element group 2377 transition  output  bypass 
    -- predecessors 2374 
    -- successors 2378 
    -- members (2) 
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xi_bbx_xnphx_xix_xi_PhiReq/phi_stmt_3757/phi_stmt_3757_sources/type_cast_3760/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xi_bbx_xnphx_xix_xi_PhiReq/phi_stmt_3757/phi_stmt_3757_sources/type_cast_3760/SplitProtocol/Update/cr
      -- 
    cp_elements(2377) <= cp_elements(2374);
    cr_19753_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2377), ack => type_cast_3760_inst_req_1); -- 
    -- CP-element group 2378 transition  input  bypass 
    -- predecessors 2377 
    -- successors 2379 
    -- members (2) 
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xi_bbx_xnphx_xix_xi_PhiReq/phi_stmt_3757/phi_stmt_3757_sources/type_cast_3760/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xi_bbx_xnphx_xix_xi_PhiReq/phi_stmt_3757/phi_stmt_3757_sources/type_cast_3760/SplitProtocol/Update/ca
      -- 
    ca_19754_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3760_inst_ack_1, ack => cp_elements(2378)); -- 
    -- CP-element group 2379 join  transition  output  bypass 
    -- predecessors 2376 2378 
    -- successors 2386 
    -- members (5) 
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xi_bbx_xnphx_xix_xi_PhiReq/phi_stmt_3757/$exit
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xi_bbx_xnphx_xix_xi_PhiReq/phi_stmt_3757/phi_stmt_3757_sources/$exit
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xi_bbx_xnphx_xix_xi_PhiReq/phi_stmt_3757/phi_stmt_3757_sources/type_cast_3760/$exit
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xi_bbx_xnphx_xix_xi_PhiReq/phi_stmt_3757/phi_stmt_3757_sources/type_cast_3760/SplitProtocol/$exit
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xi_bbx_xnphx_xix_xi_PhiReq/phi_stmt_3757/phi_stmt_3757_req
      -- 
    cp_element_group_2379: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_2379"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(2376) & cp_elements(2378);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(2379), clk => clk, reset => reset); --
    end block;
    phi_stmt_3757_req_19755_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2379), ack => phi_stmt_3757_req_0); -- 
    -- CP-element group 2380 fork  transition  bypass 
    -- predecessors 2373 
    -- successors 2381 2383 
    -- members (4) 
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xi_bbx_xnphx_xix_xi_PhiReq/phi_stmt_3764/$entry
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xi_bbx_xnphx_xix_xi_PhiReq/phi_stmt_3764/phi_stmt_3764_sources/$entry
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xi_bbx_xnphx_xix_xi_PhiReq/phi_stmt_3764/phi_stmt_3764_sources/type_cast_3767/$entry
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xi_bbx_xnphx_xix_xi_PhiReq/phi_stmt_3764/phi_stmt_3764_sources/type_cast_3767/SplitProtocol/$entry
      -- 
    cp_elements(2380) <= cp_elements(2373);
    -- CP-element group 2381 transition  output  bypass 
    -- predecessors 2380 
    -- successors 2382 
    -- members (2) 
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xi_bbx_xnphx_xix_xi_PhiReq/phi_stmt_3764/phi_stmt_3764_sources/type_cast_3767/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xi_bbx_xnphx_xix_xi_PhiReq/phi_stmt_3764/phi_stmt_3764_sources/type_cast_3767/SplitProtocol/Sample/rr
      -- 
    cp_elements(2381) <= cp_elements(2380);
    rr_19771_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2381), ack => type_cast_3767_inst_req_0); -- 
    -- CP-element group 2382 transition  input  bypass 
    -- predecessors 2381 
    -- successors 2385 
    -- members (2) 
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xi_bbx_xnphx_xix_xi_PhiReq/phi_stmt_3764/phi_stmt_3764_sources/type_cast_3767/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xi_bbx_xnphx_xix_xi_PhiReq/phi_stmt_3764/phi_stmt_3764_sources/type_cast_3767/SplitProtocol/Sample/ra
      -- 
    ra_19772_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3767_inst_ack_0, ack => cp_elements(2382)); -- 
    -- CP-element group 2383 transition  output  bypass 
    -- predecessors 2380 
    -- successors 2384 
    -- members (2) 
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xi_bbx_xnphx_xix_xi_PhiReq/phi_stmt_3764/phi_stmt_3764_sources/type_cast_3767/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xi_bbx_xnphx_xix_xi_PhiReq/phi_stmt_3764/phi_stmt_3764_sources/type_cast_3767/SplitProtocol/Update/cr
      -- 
    cp_elements(2383) <= cp_elements(2380);
    cr_19776_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2383), ack => type_cast_3767_inst_req_1); -- 
    -- CP-element group 2384 transition  input  bypass 
    -- predecessors 2383 
    -- successors 2385 
    -- members (2) 
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xi_bbx_xnphx_xix_xi_PhiReq/phi_stmt_3764/phi_stmt_3764_sources/type_cast_3767/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xi_bbx_xnphx_xix_xi_PhiReq/phi_stmt_3764/phi_stmt_3764_sources/type_cast_3767/SplitProtocol/Update/ca
      -- 
    ca_19777_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3767_inst_ack_1, ack => cp_elements(2384)); -- 
    -- CP-element group 2385 join  transition  output  bypass 
    -- predecessors 2382 2384 
    -- successors 2386 
    -- members (5) 
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xi_bbx_xnphx_xix_xi_PhiReq/phi_stmt_3764/$exit
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xi_bbx_xnphx_xix_xi_PhiReq/phi_stmt_3764/phi_stmt_3764_sources/$exit
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xi_bbx_xnphx_xix_xi_PhiReq/phi_stmt_3764/phi_stmt_3764_sources/type_cast_3767/$exit
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xi_bbx_xnphx_xix_xi_PhiReq/phi_stmt_3764/phi_stmt_3764_sources/type_cast_3767/SplitProtocol/$exit
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xi_bbx_xnphx_xix_xi_PhiReq/phi_stmt_3764/phi_stmt_3764_req
      -- 
    cp_element_group_2385: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_2385"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(2382) & cp_elements(2384);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(2385), clk => clk, reset => reset); --
    end block;
    phi_stmt_3764_req_19778_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2385), ack => phi_stmt_3764_req_0); -- 
    -- CP-element group 2386 join  transition  bypass 
    -- predecessors 2379 2385 
    -- successors 2397 
    -- members (1) 
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xi_bbx_xnphx_xix_xi_PhiReq/$exit
      -- 
    cp_element_group_2386: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_2386"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(2379) & cp_elements(2385);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(2386), clk => clk, reset => reset); --
    end block;
    -- CP-element group 2387 fork  transition  bypass 
    -- predecessors 66 
    -- successors 2388 2392 
    -- members (1) 
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xpreheader_bbx_xnphx_xix_xi_PhiReq/$entry
      -- 
    cp_elements(2387) <= cp_elements(66);
    -- CP-element group 2388 fork  transition  bypass 
    -- predecessors 2387 
    -- successors 2389 2390 
    -- members (4) 
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xpreheader_bbx_xnphx_xix_xi_PhiReq/phi_stmt_3757/$entry
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xpreheader_bbx_xnphx_xix_xi_PhiReq/phi_stmt_3757/phi_stmt_3757_sources/$entry
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xpreheader_bbx_xnphx_xix_xi_PhiReq/phi_stmt_3757/phi_stmt_3757_sources/type_cast_3760/$entry
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xpreheader_bbx_xnphx_xix_xi_PhiReq/phi_stmt_3757/phi_stmt_3757_sources/type_cast_3760/SplitProtocol/$entry
      -- 
    cp_elements(2388) <= cp_elements(2387);
    -- CP-element group 2389 transition  bypass 
    -- predecessors 2388 
    -- successors 2391 
    -- members (4) 
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xpreheader_bbx_xnphx_xix_xi_PhiReq/phi_stmt_3757/phi_stmt_3757_sources/type_cast_3760/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xpreheader_bbx_xnphx_xix_xi_PhiReq/phi_stmt_3757/phi_stmt_3757_sources/type_cast_3760/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xpreheader_bbx_xnphx_xix_xi_PhiReq/phi_stmt_3757/phi_stmt_3757_sources/type_cast_3760/SplitProtocol/Sample/rr
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xpreheader_bbx_xnphx_xix_xi_PhiReq/phi_stmt_3757/phi_stmt_3757_sources/type_cast_3760/SplitProtocol/Sample/ra
      -- 
    cp_elements(2389) <= cp_elements(2388);
    -- CP-element group 2390 transition  bypass 
    -- predecessors 2388 
    -- successors 2391 
    -- members (4) 
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xpreheader_bbx_xnphx_xix_xi_PhiReq/phi_stmt_3757/phi_stmt_3757_sources/type_cast_3760/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xpreheader_bbx_xnphx_xix_xi_PhiReq/phi_stmt_3757/phi_stmt_3757_sources/type_cast_3760/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xpreheader_bbx_xnphx_xix_xi_PhiReq/phi_stmt_3757/phi_stmt_3757_sources/type_cast_3760/SplitProtocol/Update/cr
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xpreheader_bbx_xnphx_xix_xi_PhiReq/phi_stmt_3757/phi_stmt_3757_sources/type_cast_3760/SplitProtocol/Update/ca
      -- 
    cp_elements(2390) <= cp_elements(2388);
    -- CP-element group 2391 join  transition  output  bypass 
    -- predecessors 2389 2390 
    -- successors 2396 
    -- members (5) 
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xpreheader_bbx_xnphx_xix_xi_PhiReq/phi_stmt_3757/$exit
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xpreheader_bbx_xnphx_xix_xi_PhiReq/phi_stmt_3757/phi_stmt_3757_sources/$exit
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xpreheader_bbx_xnphx_xix_xi_PhiReq/phi_stmt_3757/phi_stmt_3757_sources/type_cast_3760/$exit
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xpreheader_bbx_xnphx_xix_xi_PhiReq/phi_stmt_3757/phi_stmt_3757_sources/type_cast_3760/SplitProtocol/$exit
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xpreheader_bbx_xnphx_xix_xi_PhiReq/phi_stmt_3757/phi_stmt_3757_req
      -- 
    cp_element_group_2391: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_2391"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(2389) & cp_elements(2390);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(2391), clk => clk, reset => reset); --
    end block;
    phi_stmt_3757_req_19804_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2391), ack => phi_stmt_3757_req_1); -- 
    -- CP-element group 2392 fork  transition  bypass 
    -- predecessors 2387 
    -- successors 2393 2394 
    -- members (4) 
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xpreheader_bbx_xnphx_xix_xi_PhiReq/phi_stmt_3764/$entry
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xpreheader_bbx_xnphx_xix_xi_PhiReq/phi_stmt_3764/phi_stmt_3764_sources/$entry
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xpreheader_bbx_xnphx_xix_xi_PhiReq/phi_stmt_3764/phi_stmt_3764_sources/type_cast_3767/$entry
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xpreheader_bbx_xnphx_xix_xi_PhiReq/phi_stmt_3764/phi_stmt_3764_sources/type_cast_3767/SplitProtocol/$entry
      -- 
    cp_elements(2392) <= cp_elements(2387);
    -- CP-element group 2393 transition  bypass 
    -- predecessors 2392 
    -- successors 2395 
    -- members (4) 
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xpreheader_bbx_xnphx_xix_xi_PhiReq/phi_stmt_3764/phi_stmt_3764_sources/type_cast_3767/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xpreheader_bbx_xnphx_xix_xi_PhiReq/phi_stmt_3764/phi_stmt_3764_sources/type_cast_3767/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xpreheader_bbx_xnphx_xix_xi_PhiReq/phi_stmt_3764/phi_stmt_3764_sources/type_cast_3767/SplitProtocol/Sample/rr
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xpreheader_bbx_xnphx_xix_xi_PhiReq/phi_stmt_3764/phi_stmt_3764_sources/type_cast_3767/SplitProtocol/Sample/ra
      -- 
    cp_elements(2393) <= cp_elements(2392);
    -- CP-element group 2394 transition  bypass 
    -- predecessors 2392 
    -- successors 2395 
    -- members (4) 
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xpreheader_bbx_xnphx_xix_xi_PhiReq/phi_stmt_3764/phi_stmt_3764_sources/type_cast_3767/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xpreheader_bbx_xnphx_xix_xi_PhiReq/phi_stmt_3764/phi_stmt_3764_sources/type_cast_3767/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xpreheader_bbx_xnphx_xix_xi_PhiReq/phi_stmt_3764/phi_stmt_3764_sources/type_cast_3767/SplitProtocol/Update/cr
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xpreheader_bbx_xnphx_xix_xi_PhiReq/phi_stmt_3764/phi_stmt_3764_sources/type_cast_3767/SplitProtocol/Update/ca
      -- 
    cp_elements(2394) <= cp_elements(2392);
    -- CP-element group 2395 join  transition  output  bypass 
    -- predecessors 2393 2394 
    -- successors 2396 
    -- members (5) 
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xpreheader_bbx_xnphx_xix_xi_PhiReq/phi_stmt_3764/$exit
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xpreheader_bbx_xnphx_xix_xi_PhiReq/phi_stmt_3764/phi_stmt_3764_sources/$exit
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xpreheader_bbx_xnphx_xix_xi_PhiReq/phi_stmt_3764/phi_stmt_3764_sources/type_cast_3767/$exit
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xpreheader_bbx_xnphx_xix_xi_PhiReq/phi_stmt_3764/phi_stmt_3764_sources/type_cast_3767/SplitProtocol/$exit
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xpreheader_bbx_xnphx_xix_xi_PhiReq/phi_stmt_3764/phi_stmt_3764_req
      -- 
    cp_element_group_2395: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_2395"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(2393) & cp_elements(2394);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(2395), clk => clk, reset => reset); --
    end block;
    phi_stmt_3764_req_19827_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2395), ack => phi_stmt_3764_req_1); -- 
    -- CP-element group 2396 join  transition  bypass 
    -- predecessors 2391 2395 
    -- successors 2397 
    -- members (1) 
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xix_xpreheader_bbx_xnphx_xix_xi_PhiReq/$exit
      -- 
    cp_element_group_2396: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_2396"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(2391) & cp_elements(2395);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(2396), clk => clk, reset => reset); --
    end block;
    -- CP-element group 2397 merge  place  bypass 
    -- predecessors 2386 2396 
    -- successors 2398 
    -- members (1) 
      -- 	branch_block_stmt_2042/merge_stmt_3756_PhiReqMerge
      -- 
    cp_elements(2397) <= OrReduce(cp_elements(2386) & cp_elements(2396));
    -- CP-element group 2398 fork  transition  bypass 
    -- predecessors 2397 
    -- successors 2399 2400 
    -- members (1) 
      -- 	branch_block_stmt_2042/merge_stmt_3756_PhiAck/$entry
      -- 
    cp_elements(2398) <= cp_elements(2397);
    -- CP-element group 2399 transition  input  bypass 
    -- predecessors 2398 
    -- successors 2401 
    -- members (1) 
      -- 	branch_block_stmt_2042/merge_stmt_3756_PhiAck/phi_stmt_3757_ack
      -- 
    phi_stmt_3757_ack_19832_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_3757_ack_0, ack => cp_elements(2399)); -- 
    -- CP-element group 2400 transition  input  bypass 
    -- predecessors 2398 
    -- successors 2401 
    -- members (1) 
      -- 	branch_block_stmt_2042/merge_stmt_3756_PhiAck/phi_stmt_3764_ack
      -- 
    phi_stmt_3764_ack_19833_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_3764_ack_0, ack => cp_elements(2400)); -- 
    -- CP-element group 2401 join  transition  bypass 
    -- predecessors 2399 2400 
    -- successors 67 
    -- members (1) 
      -- 	branch_block_stmt_2042/merge_stmt_3756_PhiAck/$exit
      -- 
    cp_element_group_2401: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_2401"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(2399) & cp_elements(2400);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(2401), clk => clk, reset => reset); --
    end block;
    -- CP-element group 2402 fork  transition  bypass 
    -- predecessors 1124 
    -- successors 2403 2409 
    -- members (1) 
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xi_xx_x_crit_edgex_xix_xix_xloopexit_PhiReq/$entry
      -- 
    cp_elements(2402) <= cp_elements(1124);
    -- CP-element group 2403 fork  transition  bypass 
    -- predecessors 2402 
    -- successors 2404 2406 
    -- members (4) 
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xi_xx_x_crit_edgex_xix_xix_xloopexit_PhiReq/phi_stmt_3796/$entry
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xi_xx_x_crit_edgex_xix_xix_xloopexit_PhiReq/phi_stmt_3796/phi_stmt_3796_sources/$entry
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xi_xx_x_crit_edgex_xix_xix_xloopexit_PhiReq/phi_stmt_3796/phi_stmt_3796_sources/type_cast_3799/$entry
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xi_xx_x_crit_edgex_xix_xix_xloopexit_PhiReq/phi_stmt_3796/phi_stmt_3796_sources/type_cast_3799/SplitProtocol/$entry
      -- 
    cp_elements(2403) <= cp_elements(2402);
    -- CP-element group 2404 transition  output  bypass 
    -- predecessors 2403 
    -- successors 2405 
    -- members (2) 
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xi_xx_x_crit_edgex_xix_xix_xloopexit_PhiReq/phi_stmt_3796/phi_stmt_3796_sources/type_cast_3799/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xi_xx_x_crit_edgex_xix_xix_xloopexit_PhiReq/phi_stmt_3796/phi_stmt_3796_sources/type_cast_3799/SplitProtocol/Sample/rr
      -- 
    cp_elements(2404) <= cp_elements(2403);
    rr_19856_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2404), ack => type_cast_3799_inst_req_0); -- 
    -- CP-element group 2405 transition  input  bypass 
    -- predecessors 2404 
    -- successors 2408 
    -- members (2) 
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xi_xx_x_crit_edgex_xix_xix_xloopexit_PhiReq/phi_stmt_3796/phi_stmt_3796_sources/type_cast_3799/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xi_xx_x_crit_edgex_xix_xix_xloopexit_PhiReq/phi_stmt_3796/phi_stmt_3796_sources/type_cast_3799/SplitProtocol/Sample/ra
      -- 
    ra_19857_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3799_inst_ack_0, ack => cp_elements(2405)); -- 
    -- CP-element group 2406 transition  output  bypass 
    -- predecessors 2403 
    -- successors 2407 
    -- members (2) 
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xi_xx_x_crit_edgex_xix_xix_xloopexit_PhiReq/phi_stmt_3796/phi_stmt_3796_sources/type_cast_3799/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xi_xx_x_crit_edgex_xix_xix_xloopexit_PhiReq/phi_stmt_3796/phi_stmt_3796_sources/type_cast_3799/SplitProtocol/Update/cr
      -- 
    cp_elements(2406) <= cp_elements(2403);
    cr_19861_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2406), ack => type_cast_3799_inst_req_1); -- 
    -- CP-element group 2407 transition  input  bypass 
    -- predecessors 2406 
    -- successors 2408 
    -- members (2) 
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xi_xx_x_crit_edgex_xix_xix_xloopexit_PhiReq/phi_stmt_3796/phi_stmt_3796_sources/type_cast_3799/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xi_xx_x_crit_edgex_xix_xix_xloopexit_PhiReq/phi_stmt_3796/phi_stmt_3796_sources/type_cast_3799/SplitProtocol/Update/ca
      -- 
    ca_19862_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3799_inst_ack_1, ack => cp_elements(2407)); -- 
    -- CP-element group 2408 join  transition  output  bypass 
    -- predecessors 2405 2407 
    -- successors 2415 
    -- members (5) 
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xi_xx_x_crit_edgex_xix_xix_xloopexit_PhiReq/phi_stmt_3796/$exit
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xi_xx_x_crit_edgex_xix_xix_xloopexit_PhiReq/phi_stmt_3796/phi_stmt_3796_sources/$exit
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xi_xx_x_crit_edgex_xix_xix_xloopexit_PhiReq/phi_stmt_3796/phi_stmt_3796_sources/type_cast_3799/$exit
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xi_xx_x_crit_edgex_xix_xix_xloopexit_PhiReq/phi_stmt_3796/phi_stmt_3796_sources/type_cast_3799/SplitProtocol/$exit
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xi_xx_x_crit_edgex_xix_xix_xloopexit_PhiReq/phi_stmt_3796/phi_stmt_3796_req
      -- 
    cp_element_group_2408: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_2408"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(2405) & cp_elements(2407);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(2408), clk => clk, reset => reset); --
    end block;
    phi_stmt_3796_req_19863_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2408), ack => phi_stmt_3796_req_0); -- 
    -- CP-element group 2409 fork  transition  bypass 
    -- predecessors 2402 
    -- successors 2410 2412 
    -- members (4) 
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xi_xx_x_crit_edgex_xix_xix_xloopexit_PhiReq/phi_stmt_3800/$entry
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xi_xx_x_crit_edgex_xix_xix_xloopexit_PhiReq/phi_stmt_3800/phi_stmt_3800_sources/$entry
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xi_xx_x_crit_edgex_xix_xix_xloopexit_PhiReq/phi_stmt_3800/phi_stmt_3800_sources/type_cast_3803/$entry
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xi_xx_x_crit_edgex_xix_xix_xloopexit_PhiReq/phi_stmt_3800/phi_stmt_3800_sources/type_cast_3803/SplitProtocol/$entry
      -- 
    cp_elements(2409) <= cp_elements(2402);
    -- CP-element group 2410 transition  output  bypass 
    -- predecessors 2409 
    -- successors 2411 
    -- members (2) 
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xi_xx_x_crit_edgex_xix_xix_xloopexit_PhiReq/phi_stmt_3800/phi_stmt_3800_sources/type_cast_3803/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xi_xx_x_crit_edgex_xix_xix_xloopexit_PhiReq/phi_stmt_3800/phi_stmt_3800_sources/type_cast_3803/SplitProtocol/Sample/rr
      -- 
    cp_elements(2410) <= cp_elements(2409);
    rr_19879_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2410), ack => type_cast_3803_inst_req_0); -- 
    -- CP-element group 2411 transition  input  bypass 
    -- predecessors 2410 
    -- successors 2414 
    -- members (2) 
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xi_xx_x_crit_edgex_xix_xix_xloopexit_PhiReq/phi_stmt_3800/phi_stmt_3800_sources/type_cast_3803/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xi_xx_x_crit_edgex_xix_xix_xloopexit_PhiReq/phi_stmt_3800/phi_stmt_3800_sources/type_cast_3803/SplitProtocol/Sample/ra
      -- 
    ra_19880_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3803_inst_ack_0, ack => cp_elements(2411)); -- 
    -- CP-element group 2412 transition  output  bypass 
    -- predecessors 2409 
    -- successors 2413 
    -- members (2) 
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xi_xx_x_crit_edgex_xix_xix_xloopexit_PhiReq/phi_stmt_3800/phi_stmt_3800_sources/type_cast_3803/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xi_xx_x_crit_edgex_xix_xix_xloopexit_PhiReq/phi_stmt_3800/phi_stmt_3800_sources/type_cast_3803/SplitProtocol/Update/cr
      -- 
    cp_elements(2412) <= cp_elements(2409);
    cr_19884_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2412), ack => type_cast_3803_inst_req_1); -- 
    -- CP-element group 2413 transition  input  bypass 
    -- predecessors 2412 
    -- successors 2414 
    -- members (2) 
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xi_xx_x_crit_edgex_xix_xix_xloopexit_PhiReq/phi_stmt_3800/phi_stmt_3800_sources/type_cast_3803/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xi_xx_x_crit_edgex_xix_xix_xloopexit_PhiReq/phi_stmt_3800/phi_stmt_3800_sources/type_cast_3803/SplitProtocol/Update/ca
      -- 
    ca_19885_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3803_inst_ack_1, ack => cp_elements(2413)); -- 
    -- CP-element group 2414 join  transition  output  bypass 
    -- predecessors 2411 2413 
    -- successors 2415 
    -- members (5) 
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xi_xx_x_crit_edgex_xix_xix_xloopexit_PhiReq/phi_stmt_3800/$exit
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xi_xx_x_crit_edgex_xix_xix_xloopexit_PhiReq/phi_stmt_3800/phi_stmt_3800_sources/$exit
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xi_xx_x_crit_edgex_xix_xix_xloopexit_PhiReq/phi_stmt_3800/phi_stmt_3800_sources/type_cast_3803/$exit
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xi_xx_x_crit_edgex_xix_xix_xloopexit_PhiReq/phi_stmt_3800/phi_stmt_3800_sources/type_cast_3803/SplitProtocol/$exit
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xi_xx_x_crit_edgex_xix_xix_xloopexit_PhiReq/phi_stmt_3800/phi_stmt_3800_req
      -- 
    cp_element_group_2414: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_2414"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(2411) & cp_elements(2413);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(2414), clk => clk, reset => reset); --
    end block;
    phi_stmt_3800_req_19886_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2414), ack => phi_stmt_3800_req_0); -- 
    -- CP-element group 2415 join  transition  bypass 
    -- predecessors 2408 2414 
    -- successors 2416 
    -- members (1) 
      -- 	branch_block_stmt_2042/bbx_xnphx_xix_xi_xx_x_crit_edgex_xix_xix_xloopexit_PhiReq/$exit
      -- 
    cp_element_group_2415: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_2415"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(2408) & cp_elements(2414);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(2415), clk => clk, reset => reset); --
    end block;
    -- CP-element group 2416 place  bypass 
    -- predecessors 2415 
    -- successors 2417 
    -- members (1) 
      -- 	branch_block_stmt_2042/merge_stmt_3795_PhiReqMerge
      -- 
    cp_elements(2416) <= cp_elements(2415);
    -- CP-element group 2417 fork  transition  bypass 
    -- predecessors 2416 
    -- successors 2418 2419 
    -- members (1) 
      -- 	branch_block_stmt_2042/merge_stmt_3795_PhiAck/$entry
      -- 
    cp_elements(2417) <= cp_elements(2416);
    -- CP-element group 2418 transition  input  bypass 
    -- predecessors 2417 
    -- successors 2420 
    -- members (1) 
      -- 	branch_block_stmt_2042/merge_stmt_3795_PhiAck/phi_stmt_3796_ack
      -- 
    phi_stmt_3796_ack_19891_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_3796_ack_0, ack => cp_elements(2418)); -- 
    -- CP-element group 2419 transition  input  bypass 
    -- predecessors 2417 
    -- successors 2420 
    -- members (1) 
      -- 	branch_block_stmt_2042/merge_stmt_3795_PhiAck/phi_stmt_3800_ack
      -- 
    phi_stmt_3800_ack_19892_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_3800_ack_0, ack => cp_elements(2419)); -- 
    -- CP-element group 2420 join  transition  bypass 
    -- predecessors 2418 2419 
    -- successors 69 
    -- members (1) 
      -- 	branch_block_stmt_2042/merge_stmt_3795_PhiAck/$exit
      -- 
    cp_element_group_2420: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_2420"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(2418) & cp_elements(2419);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(2420), clk => clk, reset => reset); --
    end block;
    -- CP-element group 2421 fork  transition  bypass 
    -- predecessors 1102 
    -- successors 2422 2426 
    -- members (1) 
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xi_xx_x_crit_edgex_xix_xi_PhiReq/$entry
      -- 
    cp_elements(2421) <= cp_elements(1102);
    -- CP-element group 2422 fork  transition  bypass 
    -- predecessors 2421 
    -- successors 2423 2424 
    -- members (4) 
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xi_xx_x_crit_edgex_xix_xi_PhiReq/phi_stmt_3807/$entry
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xi_xx_x_crit_edgex_xix_xi_PhiReq/phi_stmt_3807/phi_stmt_3807_sources/$entry
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xi_xx_x_crit_edgex_xix_xi_PhiReq/phi_stmt_3807/phi_stmt_3807_sources/type_cast_3813/$entry
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xi_xx_x_crit_edgex_xix_xi_PhiReq/phi_stmt_3807/phi_stmt_3807_sources/type_cast_3813/SplitProtocol/$entry
      -- 
    cp_elements(2422) <= cp_elements(2421);
    -- CP-element group 2423 transition  bypass 
    -- predecessors 2422 
    -- successors 2425 
    -- members (4) 
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xi_xx_x_crit_edgex_xix_xi_PhiReq/phi_stmt_3807/phi_stmt_3807_sources/type_cast_3813/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xi_xx_x_crit_edgex_xix_xi_PhiReq/phi_stmt_3807/phi_stmt_3807_sources/type_cast_3813/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xi_xx_x_crit_edgex_xix_xi_PhiReq/phi_stmt_3807/phi_stmt_3807_sources/type_cast_3813/SplitProtocol/Sample/rr
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xi_xx_x_crit_edgex_xix_xi_PhiReq/phi_stmt_3807/phi_stmt_3807_sources/type_cast_3813/SplitProtocol/Sample/ra
      -- 
    cp_elements(2423) <= cp_elements(2422);
    -- CP-element group 2424 transition  bypass 
    -- predecessors 2422 
    -- successors 2425 
    -- members (4) 
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xi_xx_x_crit_edgex_xix_xi_PhiReq/phi_stmt_3807/phi_stmt_3807_sources/type_cast_3813/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xi_xx_x_crit_edgex_xix_xi_PhiReq/phi_stmt_3807/phi_stmt_3807_sources/type_cast_3813/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xi_xx_x_crit_edgex_xix_xi_PhiReq/phi_stmt_3807/phi_stmt_3807_sources/type_cast_3813/SplitProtocol/Update/cr
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xi_xx_x_crit_edgex_xix_xi_PhiReq/phi_stmt_3807/phi_stmt_3807_sources/type_cast_3813/SplitProtocol/Update/ca
      -- 
    cp_elements(2424) <= cp_elements(2422);
    -- CP-element group 2425 join  transition  output  bypass 
    -- predecessors 2423 2424 
    -- successors 2430 
    -- members (5) 
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xi_xx_x_crit_edgex_xix_xi_PhiReq/phi_stmt_3807/$exit
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xi_xx_x_crit_edgex_xix_xi_PhiReq/phi_stmt_3807/phi_stmt_3807_sources/$exit
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xi_xx_x_crit_edgex_xix_xi_PhiReq/phi_stmt_3807/phi_stmt_3807_sources/type_cast_3813/$exit
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xi_xx_x_crit_edgex_xix_xi_PhiReq/phi_stmt_3807/phi_stmt_3807_sources/type_cast_3813/SplitProtocol/$exit
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xi_xx_x_crit_edgex_xix_xi_PhiReq/phi_stmt_3807/phi_stmt_3807_req
      -- 
    cp_element_group_2425: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_2425"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(2423) & cp_elements(2424);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(2425), clk => clk, reset => reset); --
    end block;
    phi_stmt_3807_req_19918_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2425), ack => phi_stmt_3807_req_0); -- 
    -- CP-element group 2426 fork  transition  bypass 
    -- predecessors 2421 
    -- successors 2427 2428 
    -- members (4) 
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xi_xx_x_crit_edgex_xix_xi_PhiReq/phi_stmt_3814/$entry
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xi_xx_x_crit_edgex_xix_xi_PhiReq/phi_stmt_3814/phi_stmt_3814_sources/$entry
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xi_xx_x_crit_edgex_xix_xi_PhiReq/phi_stmt_3814/phi_stmt_3814_sources/type_cast_3820/$entry
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xi_xx_x_crit_edgex_xix_xi_PhiReq/phi_stmt_3814/phi_stmt_3814_sources/type_cast_3820/SplitProtocol/$entry
      -- 
    cp_elements(2426) <= cp_elements(2421);
    -- CP-element group 2427 transition  bypass 
    -- predecessors 2426 
    -- successors 2429 
    -- members (4) 
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xi_xx_x_crit_edgex_xix_xi_PhiReq/phi_stmt_3814/phi_stmt_3814_sources/type_cast_3820/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xi_xx_x_crit_edgex_xix_xi_PhiReq/phi_stmt_3814/phi_stmt_3814_sources/type_cast_3820/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xi_xx_x_crit_edgex_xix_xi_PhiReq/phi_stmt_3814/phi_stmt_3814_sources/type_cast_3820/SplitProtocol/Sample/rr
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xi_xx_x_crit_edgex_xix_xi_PhiReq/phi_stmt_3814/phi_stmt_3814_sources/type_cast_3820/SplitProtocol/Sample/ra
      -- 
    cp_elements(2427) <= cp_elements(2426);
    -- CP-element group 2428 transition  bypass 
    -- predecessors 2426 
    -- successors 2429 
    -- members (4) 
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xi_xx_x_crit_edgex_xix_xi_PhiReq/phi_stmt_3814/phi_stmt_3814_sources/type_cast_3820/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xi_xx_x_crit_edgex_xix_xi_PhiReq/phi_stmt_3814/phi_stmt_3814_sources/type_cast_3820/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xi_xx_x_crit_edgex_xix_xi_PhiReq/phi_stmt_3814/phi_stmt_3814_sources/type_cast_3820/SplitProtocol/Update/cr
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xi_xx_x_crit_edgex_xix_xi_PhiReq/phi_stmt_3814/phi_stmt_3814_sources/type_cast_3820/SplitProtocol/Update/ca
      -- 
    cp_elements(2428) <= cp_elements(2426);
    -- CP-element group 2429 join  transition  output  bypass 
    -- predecessors 2427 2428 
    -- successors 2430 
    -- members (5) 
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xi_xx_x_crit_edgex_xix_xi_PhiReq/phi_stmt_3814/$exit
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xi_xx_x_crit_edgex_xix_xi_PhiReq/phi_stmt_3814/phi_stmt_3814_sources/$exit
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xi_xx_x_crit_edgex_xix_xi_PhiReq/phi_stmt_3814/phi_stmt_3814_sources/type_cast_3820/$exit
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xi_xx_x_crit_edgex_xix_xi_PhiReq/phi_stmt_3814/phi_stmt_3814_sources/type_cast_3820/SplitProtocol/$exit
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xi_xx_x_crit_edgex_xix_xi_PhiReq/phi_stmt_3814/phi_stmt_3814_req
      -- 
    cp_element_group_2429: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_2429"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(2427) & cp_elements(2428);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(2429), clk => clk, reset => reset); --
    end block;
    phi_stmt_3814_req_19941_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2429), ack => phi_stmt_3814_req_0); -- 
    -- CP-element group 2430 join  transition  bypass 
    -- predecessors 2425 2429 
    -- successors 2445 
    -- members (1) 
      -- 	branch_block_stmt_2042/bbx_xnph7x_xix_xi_xx_x_crit_edgex_xix_xi_PhiReq/$exit
      -- 
    cp_element_group_2430: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_2430"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(2425) & cp_elements(2429);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(2430), clk => clk, reset => reset); --
    end block;
    -- CP-element group 2431 fork  transition  bypass 
    -- predecessors 69 
    -- successors 2432 2438 
    -- members (1) 
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xloopexit_xx_x_crit_edgex_xix_xi_PhiReq/$entry
      -- 
    cp_elements(2431) <= cp_elements(69);
    -- CP-element group 2432 fork  transition  bypass 
    -- predecessors 2431 
    -- successors 2433 2435 
    -- members (4) 
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xloopexit_xx_x_crit_edgex_xix_xi_PhiReq/phi_stmt_3807/$entry
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xloopexit_xx_x_crit_edgex_xix_xi_PhiReq/phi_stmt_3807/phi_stmt_3807_sources/$entry
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xloopexit_xx_x_crit_edgex_xix_xi_PhiReq/phi_stmt_3807/phi_stmt_3807_sources/type_cast_3813/$entry
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xloopexit_xx_x_crit_edgex_xix_xi_PhiReq/phi_stmt_3807/phi_stmt_3807_sources/type_cast_3813/SplitProtocol/$entry
      -- 
    cp_elements(2432) <= cp_elements(2431);
    -- CP-element group 2433 transition  output  bypass 
    -- predecessors 2432 
    -- successors 2434 
    -- members (2) 
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xloopexit_xx_x_crit_edgex_xix_xi_PhiReq/phi_stmt_3807/phi_stmt_3807_sources/type_cast_3813/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xloopexit_xx_x_crit_edgex_xix_xi_PhiReq/phi_stmt_3807/phi_stmt_3807_sources/type_cast_3813/SplitProtocol/Sample/rr
      -- 
    cp_elements(2433) <= cp_elements(2432);
    rr_19960_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2433), ack => type_cast_3813_inst_req_0); -- 
    -- CP-element group 2434 transition  input  bypass 
    -- predecessors 2433 
    -- successors 2437 
    -- members (2) 
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xloopexit_xx_x_crit_edgex_xix_xi_PhiReq/phi_stmt_3807/phi_stmt_3807_sources/type_cast_3813/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xloopexit_xx_x_crit_edgex_xix_xi_PhiReq/phi_stmt_3807/phi_stmt_3807_sources/type_cast_3813/SplitProtocol/Sample/ra
      -- 
    ra_19961_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3813_inst_ack_0, ack => cp_elements(2434)); -- 
    -- CP-element group 2435 transition  output  bypass 
    -- predecessors 2432 
    -- successors 2436 
    -- members (2) 
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xloopexit_xx_x_crit_edgex_xix_xi_PhiReq/phi_stmt_3807/phi_stmt_3807_sources/type_cast_3813/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xloopexit_xx_x_crit_edgex_xix_xi_PhiReq/phi_stmt_3807/phi_stmt_3807_sources/type_cast_3813/SplitProtocol/Update/cr
      -- 
    cp_elements(2435) <= cp_elements(2432);
    cr_19965_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2435), ack => type_cast_3813_inst_req_1); -- 
    -- CP-element group 2436 transition  input  bypass 
    -- predecessors 2435 
    -- successors 2437 
    -- members (2) 
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xloopexit_xx_x_crit_edgex_xix_xi_PhiReq/phi_stmt_3807/phi_stmt_3807_sources/type_cast_3813/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xloopexit_xx_x_crit_edgex_xix_xi_PhiReq/phi_stmt_3807/phi_stmt_3807_sources/type_cast_3813/SplitProtocol/Update/ca
      -- 
    ca_19966_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3813_inst_ack_1, ack => cp_elements(2436)); -- 
    -- CP-element group 2437 join  transition  output  bypass 
    -- predecessors 2434 2436 
    -- successors 2444 
    -- members (5) 
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xloopexit_xx_x_crit_edgex_xix_xi_PhiReq/phi_stmt_3807/$exit
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xloopexit_xx_x_crit_edgex_xix_xi_PhiReq/phi_stmt_3807/phi_stmt_3807_sources/$exit
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xloopexit_xx_x_crit_edgex_xix_xi_PhiReq/phi_stmt_3807/phi_stmt_3807_sources/type_cast_3813/$exit
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xloopexit_xx_x_crit_edgex_xix_xi_PhiReq/phi_stmt_3807/phi_stmt_3807_sources/type_cast_3813/SplitProtocol/$exit
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xloopexit_xx_x_crit_edgex_xix_xi_PhiReq/phi_stmt_3807/phi_stmt_3807_req
      -- 
    cp_element_group_2437: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_2437"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(2434) & cp_elements(2436);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(2437), clk => clk, reset => reset); --
    end block;
    phi_stmt_3807_req_19967_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2437), ack => phi_stmt_3807_req_1); -- 
    -- CP-element group 2438 fork  transition  bypass 
    -- predecessors 2431 
    -- successors 2439 2441 
    -- members (4) 
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xloopexit_xx_x_crit_edgex_xix_xi_PhiReq/phi_stmt_3814/$entry
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xloopexit_xx_x_crit_edgex_xix_xi_PhiReq/phi_stmt_3814/phi_stmt_3814_sources/$entry
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xloopexit_xx_x_crit_edgex_xix_xi_PhiReq/phi_stmt_3814/phi_stmt_3814_sources/type_cast_3820/$entry
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xloopexit_xx_x_crit_edgex_xix_xi_PhiReq/phi_stmt_3814/phi_stmt_3814_sources/type_cast_3820/SplitProtocol/$entry
      -- 
    cp_elements(2438) <= cp_elements(2431);
    -- CP-element group 2439 transition  output  bypass 
    -- predecessors 2438 
    -- successors 2440 
    -- members (2) 
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xloopexit_xx_x_crit_edgex_xix_xi_PhiReq/phi_stmt_3814/phi_stmt_3814_sources/type_cast_3820/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xloopexit_xx_x_crit_edgex_xix_xi_PhiReq/phi_stmt_3814/phi_stmt_3814_sources/type_cast_3820/SplitProtocol/Sample/rr
      -- 
    cp_elements(2439) <= cp_elements(2438);
    rr_19983_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2439), ack => type_cast_3820_inst_req_0); -- 
    -- CP-element group 2440 transition  input  bypass 
    -- predecessors 2439 
    -- successors 2443 
    -- members (2) 
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xloopexit_xx_x_crit_edgex_xix_xi_PhiReq/phi_stmt_3814/phi_stmt_3814_sources/type_cast_3820/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xloopexit_xx_x_crit_edgex_xix_xi_PhiReq/phi_stmt_3814/phi_stmt_3814_sources/type_cast_3820/SplitProtocol/Sample/ra
      -- 
    ra_19984_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3820_inst_ack_0, ack => cp_elements(2440)); -- 
    -- CP-element group 2441 transition  output  bypass 
    -- predecessors 2438 
    -- successors 2442 
    -- members (2) 
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xloopexit_xx_x_crit_edgex_xix_xi_PhiReq/phi_stmt_3814/phi_stmt_3814_sources/type_cast_3820/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xloopexit_xx_x_crit_edgex_xix_xi_PhiReq/phi_stmt_3814/phi_stmt_3814_sources/type_cast_3820/SplitProtocol/Update/cr
      -- 
    cp_elements(2441) <= cp_elements(2438);
    cr_19988_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2441), ack => type_cast_3820_inst_req_1); -- 
    -- CP-element group 2442 transition  input  bypass 
    -- predecessors 2441 
    -- successors 2443 
    -- members (2) 
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xloopexit_xx_x_crit_edgex_xix_xi_PhiReq/phi_stmt_3814/phi_stmt_3814_sources/type_cast_3820/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xloopexit_xx_x_crit_edgex_xix_xi_PhiReq/phi_stmt_3814/phi_stmt_3814_sources/type_cast_3820/SplitProtocol/Update/ca
      -- 
    ca_19989_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3820_inst_ack_1, ack => cp_elements(2442)); -- 
    -- CP-element group 2443 join  transition  output  bypass 
    -- predecessors 2440 2442 
    -- successors 2444 
    -- members (5) 
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xloopexit_xx_x_crit_edgex_xix_xi_PhiReq/phi_stmt_3814/$exit
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xloopexit_xx_x_crit_edgex_xix_xi_PhiReq/phi_stmt_3814/phi_stmt_3814_sources/$exit
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xloopexit_xx_x_crit_edgex_xix_xi_PhiReq/phi_stmt_3814/phi_stmt_3814_sources/type_cast_3820/$exit
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xloopexit_xx_x_crit_edgex_xix_xi_PhiReq/phi_stmt_3814/phi_stmt_3814_sources/type_cast_3820/SplitProtocol/$exit
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xloopexit_xx_x_crit_edgex_xix_xi_PhiReq/phi_stmt_3814/phi_stmt_3814_req
      -- 
    cp_element_group_2443: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_2443"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(2440) & cp_elements(2442);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(2443), clk => clk, reset => reset); --
    end block;
    phi_stmt_3814_req_19990_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2443), ack => phi_stmt_3814_req_1); -- 
    -- CP-element group 2444 join  transition  bypass 
    -- predecessors 2437 2443 
    -- successors 2445 
    -- members (1) 
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xix_xloopexit_xx_x_crit_edgex_xix_xi_PhiReq/$exit
      -- 
    cp_element_group_2444: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_2444"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(2437) & cp_elements(2443);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(2444), clk => clk, reset => reset); --
    end block;
    -- CP-element group 2445 merge  place  bypass 
    -- predecessors 2430 2444 
    -- successors 2446 
    -- members (1) 
      -- 	branch_block_stmt_2042/merge_stmt_3806_PhiReqMerge
      -- 
    cp_elements(2445) <= OrReduce(cp_elements(2430) & cp_elements(2444));
    -- CP-element group 2446 fork  transition  bypass 
    -- predecessors 2445 
    -- successors 2447 2448 
    -- members (1) 
      -- 	branch_block_stmt_2042/merge_stmt_3806_PhiAck/$entry
      -- 
    cp_elements(2446) <= cp_elements(2445);
    -- CP-element group 2447 transition  input  bypass 
    -- predecessors 2446 
    -- successors 2449 
    -- members (1) 
      -- 	branch_block_stmt_2042/merge_stmt_3806_PhiAck/phi_stmt_3807_ack
      -- 
    phi_stmt_3807_ack_19995_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_3807_ack_0, ack => cp_elements(2447)); -- 
    -- CP-element group 2448 transition  input  bypass 
    -- predecessors 2446 
    -- successors 2449 
    -- members (1) 
      -- 	branch_block_stmt_2042/merge_stmt_3806_PhiAck/phi_stmt_3814_ack
      -- 
    phi_stmt_3814_ack_19996_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_3814_ack_0, ack => cp_elements(2448)); -- 
    -- CP-element group 2449 join  transition  bypass 
    -- predecessors 2447 2448 
    -- successors 70 
    -- members (1) 
      -- 	branch_block_stmt_2042/merge_stmt_3806_PhiAck/$exit
      -- 
    cp_element_group_2449: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_2449"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(2447) & cp_elements(2448);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(2449), clk => clk, reset => reset); --
    end block;
    -- CP-element group 2450 transition  output  bypass 
    -- predecessors 1146 
    -- successors 2451 
    -- members (2) 
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xi_udiv32x_xexitx_xpreheaderx_xi_PhiReq/phi_stmt_3845/phi_stmt_3845_sources/type_cast_3848/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xi_udiv32x_xexitx_xpreheaderx_xi_PhiReq/phi_stmt_3845/phi_stmt_3845_sources/type_cast_3848/SplitProtocol/Sample/rr
      -- 
    cp_elements(2450) <= cp_elements(1146);
    rr_20019_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2450), ack => type_cast_3848_inst_req_0); -- 
    -- CP-element group 2451 transition  input  bypass 
    -- predecessors 2450 
    -- successors 2454 
    -- members (2) 
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xi_udiv32x_xexitx_xpreheaderx_xi_PhiReq/phi_stmt_3845/phi_stmt_3845_sources/type_cast_3848/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xi_udiv32x_xexitx_xpreheaderx_xi_PhiReq/phi_stmt_3845/phi_stmt_3845_sources/type_cast_3848/SplitProtocol/Sample/ra
      -- 
    ra_20020_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3848_inst_ack_0, ack => cp_elements(2451)); -- 
    -- CP-element group 2452 transition  output  bypass 
    -- predecessors 1146 
    -- successors 2453 
    -- members (2) 
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xi_udiv32x_xexitx_xpreheaderx_xi_PhiReq/phi_stmt_3845/phi_stmt_3845_sources/type_cast_3848/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xi_udiv32x_xexitx_xpreheaderx_xi_PhiReq/phi_stmt_3845/phi_stmt_3845_sources/type_cast_3848/SplitProtocol/Update/cr
      -- 
    cp_elements(2452) <= cp_elements(1146);
    cr_20024_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2452), ack => type_cast_3848_inst_req_1); -- 
    -- CP-element group 2453 transition  input  bypass 
    -- predecessors 2452 
    -- successors 2454 
    -- members (2) 
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xi_udiv32x_xexitx_xpreheaderx_xi_PhiReq/phi_stmt_3845/phi_stmt_3845_sources/type_cast_3848/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xi_udiv32x_xexitx_xpreheaderx_xi_PhiReq/phi_stmt_3845/phi_stmt_3845_sources/type_cast_3848/SplitProtocol/Update/ca
      -- 
    ca_20025_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3848_inst_ack_1, ack => cp_elements(2453)); -- 
    -- CP-element group 2454 join  transition  place  output  bypass 
    -- predecessors 2451 2453 
    -- successors 2455 
    -- members (8) 
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xi_udiv32x_xexitx_xpreheaderx_xi_PhiReq/$exit
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xi_udiv32x_xexitx_xpreheaderx_xi_PhiReq/phi_stmt_3845/$exit
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xi_udiv32x_xexitx_xpreheaderx_xi_PhiReq/phi_stmt_3845/phi_stmt_3845_sources/$exit
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xi_udiv32x_xexitx_xpreheaderx_xi_PhiReq/phi_stmt_3845/phi_stmt_3845_sources/type_cast_3848/$exit
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xi_udiv32x_xexitx_xpreheaderx_xi_PhiReq/phi_stmt_3845/phi_stmt_3845_sources/type_cast_3848/SplitProtocol/$exit
      -- 	branch_block_stmt_2042/xx_x_crit_edgex_xix_xi_udiv32x_xexitx_xpreheaderx_xi_PhiReq/phi_stmt_3845/phi_stmt_3845_req
      -- 	branch_block_stmt_2042/merge_stmt_3844_PhiReqMerge
      -- 	branch_block_stmt_2042/merge_stmt_3844_PhiAck/$entry
      -- 
    cp_element_group_2454: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_2454"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(2451) & cp_elements(2453);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(2454), clk => clk, reset => reset); --
    end block;
    phi_stmt_3845_req_20026_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2454), ack => phi_stmt_3845_req_0); -- 
    -- CP-element group 2455 transition  input  bypass 
    -- predecessors 2454 
    -- successors 72 
    -- members (2) 
      -- 	branch_block_stmt_2042/merge_stmt_3844_PhiAck/$exit
      -- 	branch_block_stmt_2042/merge_stmt_3844_PhiAck/phi_stmt_3845_ack
      -- 
    phi_stmt_3845_ack_20031_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_3845_ack_0, ack => cp_elements(2455)); -- 
    -- CP-element group 2456 fork  transition  bypass 
    -- predecessors 1220 
    -- successors 2457 2463 
    -- members (1) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xi_udiv32x_xexitx_xi_PhiReq/$entry
      -- 
    cp_elements(2456) <= cp_elements(1220);
    -- CP-element group 2457 fork  transition  bypass 
    -- predecessors 2456 
    -- successors 2458 2460 
    -- members (4) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xi_udiv32x_xexitx_xi_PhiReq/phi_stmt_3908/$entry
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xi_udiv32x_xexitx_xi_PhiReq/phi_stmt_3908/phi_stmt_3908_sources/$entry
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xi_udiv32x_xexitx_xi_PhiReq/phi_stmt_3908/phi_stmt_3908_sources/type_cast_3911/$entry
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xi_udiv32x_xexitx_xi_PhiReq/phi_stmt_3908/phi_stmt_3908_sources/type_cast_3911/SplitProtocol/$entry
      -- 
    cp_elements(2457) <= cp_elements(2456);
    -- CP-element group 2458 transition  output  bypass 
    -- predecessors 2457 
    -- successors 2459 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xi_udiv32x_xexitx_xi_PhiReq/phi_stmt_3908/phi_stmt_3908_sources/type_cast_3911/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xi_udiv32x_xexitx_xi_PhiReq/phi_stmt_3908/phi_stmt_3908_sources/type_cast_3911/SplitProtocol/Sample/rr
      -- 
    cp_elements(2458) <= cp_elements(2457);
    rr_20062_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2458), ack => type_cast_3911_inst_req_0); -- 
    -- CP-element group 2459 transition  input  bypass 
    -- predecessors 2458 
    -- successors 2462 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xi_udiv32x_xexitx_xi_PhiReq/phi_stmt_3908/phi_stmt_3908_sources/type_cast_3911/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xi_udiv32x_xexitx_xi_PhiReq/phi_stmt_3908/phi_stmt_3908_sources/type_cast_3911/SplitProtocol/Sample/ra
      -- 
    ra_20063_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3911_inst_ack_0, ack => cp_elements(2459)); -- 
    -- CP-element group 2460 transition  output  bypass 
    -- predecessors 2457 
    -- successors 2461 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xi_udiv32x_xexitx_xi_PhiReq/phi_stmt_3908/phi_stmt_3908_sources/type_cast_3911/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xi_udiv32x_xexitx_xi_PhiReq/phi_stmt_3908/phi_stmt_3908_sources/type_cast_3911/SplitProtocol/Update/cr
      -- 
    cp_elements(2460) <= cp_elements(2457);
    cr_20067_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2460), ack => type_cast_3911_inst_req_1); -- 
    -- CP-element group 2461 transition  input  bypass 
    -- predecessors 2460 
    -- successors 2462 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xi_udiv32x_xexitx_xi_PhiReq/phi_stmt_3908/phi_stmt_3908_sources/type_cast_3911/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xi_udiv32x_xexitx_xi_PhiReq/phi_stmt_3908/phi_stmt_3908_sources/type_cast_3911/SplitProtocol/Update/ca
      -- 
    ca_20068_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3911_inst_ack_1, ack => cp_elements(2461)); -- 
    -- CP-element group 2462 join  transition  output  bypass 
    -- predecessors 2459 2461 
    -- successors 2475 
    -- members (5) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xi_udiv32x_xexitx_xi_PhiReq/phi_stmt_3908/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xi_udiv32x_xexitx_xi_PhiReq/phi_stmt_3908/phi_stmt_3908_sources/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xi_udiv32x_xexitx_xi_PhiReq/phi_stmt_3908/phi_stmt_3908_sources/type_cast_3911/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xi_udiv32x_xexitx_xi_PhiReq/phi_stmt_3908/phi_stmt_3908_sources/type_cast_3911/SplitProtocol/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xi_udiv32x_xexitx_xi_PhiReq/phi_stmt_3908/phi_stmt_3908_req
      -- 
    cp_element_group_2462: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_2462"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(2459) & cp_elements(2461);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(2462), clk => clk, reset => reset); --
    end block;
    phi_stmt_3908_req_20069_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2462), ack => phi_stmt_3908_req_0); -- 
    -- CP-element group 2463 fork  transition  bypass 
    -- predecessors 2456 
    -- successors 2464 2470 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xi_udiv32x_xexitx_xi_PhiReq/phi_stmt_3915/$entry
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xi_udiv32x_xexitx_xi_PhiReq/phi_stmt_3915/phi_stmt_3915_sources/$entry
      -- 
    cp_elements(2463) <= cp_elements(2456);
    -- CP-element group 2464 fork  transition  bypass 
    -- predecessors 2463 
    -- successors 2465 2467 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xi_udiv32x_xexitx_xi_PhiReq/phi_stmt_3915/phi_stmt_3915_sources/type_cast_3918/$entry
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xi_udiv32x_xexitx_xi_PhiReq/phi_stmt_3915/phi_stmt_3915_sources/type_cast_3918/SplitProtocol/$entry
      -- 
    cp_elements(2464) <= cp_elements(2463);
    -- CP-element group 2465 transition  output  bypass 
    -- predecessors 2464 
    -- successors 2466 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xi_udiv32x_xexitx_xi_PhiReq/phi_stmt_3915/phi_stmt_3915_sources/type_cast_3918/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xi_udiv32x_xexitx_xi_PhiReq/phi_stmt_3915/phi_stmt_3915_sources/type_cast_3918/SplitProtocol/Sample/rr
      -- 
    cp_elements(2465) <= cp_elements(2464);
    rr_20085_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2465), ack => type_cast_3918_inst_req_0); -- 
    -- CP-element group 2466 transition  input  bypass 
    -- predecessors 2465 
    -- successors 2469 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xi_udiv32x_xexitx_xi_PhiReq/phi_stmt_3915/phi_stmt_3915_sources/type_cast_3918/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xi_udiv32x_xexitx_xi_PhiReq/phi_stmt_3915/phi_stmt_3915_sources/type_cast_3918/SplitProtocol/Sample/ra
      -- 
    ra_20086_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3918_inst_ack_0, ack => cp_elements(2466)); -- 
    -- CP-element group 2467 transition  output  bypass 
    -- predecessors 2464 
    -- successors 2468 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xi_udiv32x_xexitx_xi_PhiReq/phi_stmt_3915/phi_stmt_3915_sources/type_cast_3918/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xi_udiv32x_xexitx_xi_PhiReq/phi_stmt_3915/phi_stmt_3915_sources/type_cast_3918/SplitProtocol/Update/cr
      -- 
    cp_elements(2467) <= cp_elements(2464);
    cr_20090_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2467), ack => type_cast_3918_inst_req_1); -- 
    -- CP-element group 2468 transition  input  bypass 
    -- predecessors 2467 
    -- successors 2469 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xi_udiv32x_xexitx_xi_PhiReq/phi_stmt_3915/phi_stmt_3915_sources/type_cast_3918/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xi_udiv32x_xexitx_xi_PhiReq/phi_stmt_3915/phi_stmt_3915_sources/type_cast_3918/SplitProtocol/Update/ca
      -- 
    ca_20091_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3918_inst_ack_1, ack => cp_elements(2468)); -- 
    -- CP-element group 2469 join  transition  bypass 
    -- predecessors 2466 2468 
    -- successors 2474 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xi_udiv32x_xexitx_xi_PhiReq/phi_stmt_3915/phi_stmt_3915_sources/type_cast_3918/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xi_udiv32x_xexitx_xi_PhiReq/phi_stmt_3915/phi_stmt_3915_sources/type_cast_3918/SplitProtocol/$exit
      -- 
    cp_element_group_2469: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_2469"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(2466) & cp_elements(2468);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(2469), clk => clk, reset => reset); --
    end block;
    -- CP-element group 2470 fork  transition  bypass 
    -- predecessors 2463 
    -- successors 2471 2472 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xi_udiv32x_xexitx_xi_PhiReq/phi_stmt_3915/phi_stmt_3915_sources/type_cast_3920/$entry
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xi_udiv32x_xexitx_xi_PhiReq/phi_stmt_3915/phi_stmt_3915_sources/type_cast_3920/SplitProtocol/$entry
      -- 
    cp_elements(2470) <= cp_elements(2463);
    -- CP-element group 2471 transition  bypass 
    -- predecessors 2470 
    -- successors 2473 
    -- members (4) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xi_udiv32x_xexitx_xi_PhiReq/phi_stmt_3915/phi_stmt_3915_sources/type_cast_3920/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xi_udiv32x_xexitx_xi_PhiReq/phi_stmt_3915/phi_stmt_3915_sources/type_cast_3920/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xi_udiv32x_xexitx_xi_PhiReq/phi_stmt_3915/phi_stmt_3915_sources/type_cast_3920/SplitProtocol/Sample/rr
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xi_udiv32x_xexitx_xi_PhiReq/phi_stmt_3915/phi_stmt_3915_sources/type_cast_3920/SplitProtocol/Sample/ra
      -- 
    cp_elements(2471) <= cp_elements(2470);
    -- CP-element group 2472 transition  bypass 
    -- predecessors 2470 
    -- successors 2473 
    -- members (4) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xi_udiv32x_xexitx_xi_PhiReq/phi_stmt_3915/phi_stmt_3915_sources/type_cast_3920/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xi_udiv32x_xexitx_xi_PhiReq/phi_stmt_3915/phi_stmt_3915_sources/type_cast_3920/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xi_udiv32x_xexitx_xi_PhiReq/phi_stmt_3915/phi_stmt_3915_sources/type_cast_3920/SplitProtocol/Update/cr
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xi_udiv32x_xexitx_xi_PhiReq/phi_stmt_3915/phi_stmt_3915_sources/type_cast_3920/SplitProtocol/Update/ca
      -- 
    cp_elements(2472) <= cp_elements(2470);
    -- CP-element group 2473 join  transition  bypass 
    -- predecessors 2471 2472 
    -- successors 2474 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xi_udiv32x_xexitx_xi_PhiReq/phi_stmt_3915/phi_stmt_3915_sources/type_cast_3920/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xi_udiv32x_xexitx_xi_PhiReq/phi_stmt_3915/phi_stmt_3915_sources/type_cast_3920/SplitProtocol/$exit
      -- 
    cp_element_group_2473: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_2473"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(2471) & cp_elements(2472);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(2473), clk => clk, reset => reset); --
    end block;
    -- CP-element group 2474 join  transition  output  bypass 
    -- predecessors 2469 2473 
    -- successors 2475 
    -- members (3) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xi_udiv32x_xexitx_xi_PhiReq/phi_stmt_3915/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xi_udiv32x_xexitx_xi_PhiReq/phi_stmt_3915/phi_stmt_3915_sources/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xi_udiv32x_xexitx_xi_PhiReq/phi_stmt_3915/phi_stmt_3915_req
      -- 
    cp_element_group_2474: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_2474"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(2469) & cp_elements(2473);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(2474), clk => clk, reset => reset); --
    end block;
    phi_stmt_3915_req_20108_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2474), ack => phi_stmt_3915_req_0); -- 
    -- CP-element group 2475 join  transition  bypass 
    -- predecessors 2462 2474 
    -- successors 2494 
    -- members (1) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xi_udiv32x_xexitx_xi_PhiReq/$exit
      -- 
    cp_element_group_2475: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_2475"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(2462) & cp_elements(2474);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(2475), clk => clk, reset => reset); --
    end block;
    -- CP-element group 2476 fork  transition  bypass 
    -- predecessors 74 
    -- successors 2477 2481 
    -- members (1) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xpreheader_udiv32x_xexitx_xi_PhiReq/$entry
      -- 
    cp_elements(2476) <= cp_elements(74);
    -- CP-element group 2477 fork  transition  bypass 
    -- predecessors 2476 
    -- successors 2478 2479 
    -- members (4) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xpreheader_udiv32x_xexitx_xi_PhiReq/phi_stmt_3908/$entry
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xpreheader_udiv32x_xexitx_xi_PhiReq/phi_stmt_3908/phi_stmt_3908_sources/$entry
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xpreheader_udiv32x_xexitx_xi_PhiReq/phi_stmt_3908/phi_stmt_3908_sources/type_cast_3911/$entry
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xpreheader_udiv32x_xexitx_xi_PhiReq/phi_stmt_3908/phi_stmt_3908_sources/type_cast_3911/SplitProtocol/$entry
      -- 
    cp_elements(2477) <= cp_elements(2476);
    -- CP-element group 2478 transition  bypass 
    -- predecessors 2477 
    -- successors 2480 
    -- members (4) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xpreheader_udiv32x_xexitx_xi_PhiReq/phi_stmt_3908/phi_stmt_3908_sources/type_cast_3911/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xpreheader_udiv32x_xexitx_xi_PhiReq/phi_stmt_3908/phi_stmt_3908_sources/type_cast_3911/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xpreheader_udiv32x_xexitx_xi_PhiReq/phi_stmt_3908/phi_stmt_3908_sources/type_cast_3911/SplitProtocol/Sample/rr
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xpreheader_udiv32x_xexitx_xi_PhiReq/phi_stmt_3908/phi_stmt_3908_sources/type_cast_3911/SplitProtocol/Sample/ra
      -- 
    cp_elements(2478) <= cp_elements(2477);
    -- CP-element group 2479 transition  bypass 
    -- predecessors 2477 
    -- successors 2480 
    -- members (4) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xpreheader_udiv32x_xexitx_xi_PhiReq/phi_stmt_3908/phi_stmt_3908_sources/type_cast_3911/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xpreheader_udiv32x_xexitx_xi_PhiReq/phi_stmt_3908/phi_stmt_3908_sources/type_cast_3911/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xpreheader_udiv32x_xexitx_xi_PhiReq/phi_stmt_3908/phi_stmt_3908_sources/type_cast_3911/SplitProtocol/Update/cr
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xpreheader_udiv32x_xexitx_xi_PhiReq/phi_stmt_3908/phi_stmt_3908_sources/type_cast_3911/SplitProtocol/Update/ca
      -- 
    cp_elements(2479) <= cp_elements(2477);
    -- CP-element group 2480 join  transition  output  bypass 
    -- predecessors 2478 2479 
    -- successors 2493 
    -- members (5) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xpreheader_udiv32x_xexitx_xi_PhiReq/phi_stmt_3908/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xpreheader_udiv32x_xexitx_xi_PhiReq/phi_stmt_3908/phi_stmt_3908_sources/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xpreheader_udiv32x_xexitx_xi_PhiReq/phi_stmt_3908/phi_stmt_3908_sources/type_cast_3911/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xpreheader_udiv32x_xexitx_xi_PhiReq/phi_stmt_3908/phi_stmt_3908_sources/type_cast_3911/SplitProtocol/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xpreheader_udiv32x_xexitx_xi_PhiReq/phi_stmt_3908/phi_stmt_3908_req
      -- 
    cp_element_group_2480: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_2480"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(2478) & cp_elements(2479);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(2480), clk => clk, reset => reset); --
    end block;
    phi_stmt_3908_req_20134_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2480), ack => phi_stmt_3908_req_1); -- 
    -- CP-element group 2481 fork  transition  bypass 
    -- predecessors 2476 
    -- successors 2482 2486 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xpreheader_udiv32x_xexitx_xi_PhiReq/phi_stmt_3915/$entry
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xpreheader_udiv32x_xexitx_xi_PhiReq/phi_stmt_3915/phi_stmt_3915_sources/$entry
      -- 
    cp_elements(2481) <= cp_elements(2476);
    -- CP-element group 2482 fork  transition  bypass 
    -- predecessors 2481 
    -- successors 2483 2484 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xpreheader_udiv32x_xexitx_xi_PhiReq/phi_stmt_3915/phi_stmt_3915_sources/type_cast_3918/$entry
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xpreheader_udiv32x_xexitx_xi_PhiReq/phi_stmt_3915/phi_stmt_3915_sources/type_cast_3918/SplitProtocol/$entry
      -- 
    cp_elements(2482) <= cp_elements(2481);
    -- CP-element group 2483 transition  bypass 
    -- predecessors 2482 
    -- successors 2485 
    -- members (4) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xpreheader_udiv32x_xexitx_xi_PhiReq/phi_stmt_3915/phi_stmt_3915_sources/type_cast_3918/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xpreheader_udiv32x_xexitx_xi_PhiReq/phi_stmt_3915/phi_stmt_3915_sources/type_cast_3918/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xpreheader_udiv32x_xexitx_xi_PhiReq/phi_stmt_3915/phi_stmt_3915_sources/type_cast_3918/SplitProtocol/Sample/rr
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xpreheader_udiv32x_xexitx_xi_PhiReq/phi_stmt_3915/phi_stmt_3915_sources/type_cast_3918/SplitProtocol/Sample/ra
      -- 
    cp_elements(2483) <= cp_elements(2482);
    -- CP-element group 2484 transition  bypass 
    -- predecessors 2482 
    -- successors 2485 
    -- members (4) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xpreheader_udiv32x_xexitx_xi_PhiReq/phi_stmt_3915/phi_stmt_3915_sources/type_cast_3918/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xpreheader_udiv32x_xexitx_xi_PhiReq/phi_stmt_3915/phi_stmt_3915_sources/type_cast_3918/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xpreheader_udiv32x_xexitx_xi_PhiReq/phi_stmt_3915/phi_stmt_3915_sources/type_cast_3918/SplitProtocol/Update/cr
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xpreheader_udiv32x_xexitx_xi_PhiReq/phi_stmt_3915/phi_stmt_3915_sources/type_cast_3918/SplitProtocol/Update/ca
      -- 
    cp_elements(2484) <= cp_elements(2482);
    -- CP-element group 2485 join  transition  bypass 
    -- predecessors 2483 2484 
    -- successors 2492 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xpreheader_udiv32x_xexitx_xi_PhiReq/phi_stmt_3915/phi_stmt_3915_sources/type_cast_3918/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xpreheader_udiv32x_xexitx_xi_PhiReq/phi_stmt_3915/phi_stmt_3915_sources/type_cast_3918/SplitProtocol/$exit
      -- 
    cp_element_group_2485: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_2485"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(2483) & cp_elements(2484);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(2485), clk => clk, reset => reset); --
    end block;
    -- CP-element group 2486 fork  transition  bypass 
    -- predecessors 2481 
    -- successors 2487 2489 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xpreheader_udiv32x_xexitx_xi_PhiReq/phi_stmt_3915/phi_stmt_3915_sources/type_cast_3920/$entry
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xpreheader_udiv32x_xexitx_xi_PhiReq/phi_stmt_3915/phi_stmt_3915_sources/type_cast_3920/SplitProtocol/$entry
      -- 
    cp_elements(2486) <= cp_elements(2481);
    -- CP-element group 2487 transition  output  bypass 
    -- predecessors 2486 
    -- successors 2488 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xpreheader_udiv32x_xexitx_xi_PhiReq/phi_stmt_3915/phi_stmt_3915_sources/type_cast_3920/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xpreheader_udiv32x_xexitx_xi_PhiReq/phi_stmt_3915/phi_stmt_3915_sources/type_cast_3920/SplitProtocol/Sample/rr
      -- 
    cp_elements(2487) <= cp_elements(2486);
    rr_20166_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2487), ack => type_cast_3920_inst_req_0); -- 
    -- CP-element group 2488 transition  input  bypass 
    -- predecessors 2487 
    -- successors 2491 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xpreheader_udiv32x_xexitx_xi_PhiReq/phi_stmt_3915/phi_stmt_3915_sources/type_cast_3920/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xpreheader_udiv32x_xexitx_xi_PhiReq/phi_stmt_3915/phi_stmt_3915_sources/type_cast_3920/SplitProtocol/Sample/ra
      -- 
    ra_20167_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3920_inst_ack_0, ack => cp_elements(2488)); -- 
    -- CP-element group 2489 transition  output  bypass 
    -- predecessors 2486 
    -- successors 2490 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xpreheader_udiv32x_xexitx_xi_PhiReq/phi_stmt_3915/phi_stmt_3915_sources/type_cast_3920/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xpreheader_udiv32x_xexitx_xi_PhiReq/phi_stmt_3915/phi_stmt_3915_sources/type_cast_3920/SplitProtocol/Update/cr
      -- 
    cp_elements(2489) <= cp_elements(2486);
    cr_20171_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2489), ack => type_cast_3920_inst_req_1); -- 
    -- CP-element group 2490 transition  input  bypass 
    -- predecessors 2489 
    -- successors 2491 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xpreheader_udiv32x_xexitx_xi_PhiReq/phi_stmt_3915/phi_stmt_3915_sources/type_cast_3920/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xpreheader_udiv32x_xexitx_xi_PhiReq/phi_stmt_3915/phi_stmt_3915_sources/type_cast_3920/SplitProtocol/Update/ca
      -- 
    ca_20172_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3920_inst_ack_1, ack => cp_elements(2490)); -- 
    -- CP-element group 2491 join  transition  bypass 
    -- predecessors 2488 2490 
    -- successors 2492 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xpreheader_udiv32x_xexitx_xi_PhiReq/phi_stmt_3915/phi_stmt_3915_sources/type_cast_3920/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xpreheader_udiv32x_xexitx_xi_PhiReq/phi_stmt_3915/phi_stmt_3915_sources/type_cast_3920/SplitProtocol/$exit
      -- 
    cp_element_group_2491: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_2491"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(2488) & cp_elements(2490);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(2491), clk => clk, reset => reset); --
    end block;
    -- CP-element group 2492 join  transition  output  bypass 
    -- predecessors 2485 2491 
    -- successors 2493 
    -- members (3) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xpreheader_udiv32x_xexitx_xi_PhiReq/phi_stmt_3915/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xpreheader_udiv32x_xexitx_xi_PhiReq/phi_stmt_3915/phi_stmt_3915_sources/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xpreheader_udiv32x_xexitx_xi_PhiReq/phi_stmt_3915/phi_stmt_3915_req
      -- 
    cp_element_group_2492: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_2492"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(2485) & cp_elements(2491);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(2492), clk => clk, reset => reset); --
    end block;
    phi_stmt_3915_req_20173_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2492), ack => phi_stmt_3915_req_1); -- 
    -- CP-element group 2493 join  transition  bypass 
    -- predecessors 2480 2492 
    -- successors 2494 
    -- members (1) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xix_xpreheader_udiv32x_xexitx_xi_PhiReq/$exit
      -- 
    cp_element_group_2493: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_2493"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(2480) & cp_elements(2492);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(2493), clk => clk, reset => reset); --
    end block;
    -- CP-element group 2494 merge  place  bypass 
    -- predecessors 2475 2493 
    -- successors 2495 
    -- members (1) 
      -- 	branch_block_stmt_2042/merge_stmt_3907_PhiReqMerge
      -- 
    cp_elements(2494) <= OrReduce(cp_elements(2475) & cp_elements(2493));
    -- CP-element group 2495 fork  transition  bypass 
    -- predecessors 2494 
    -- successors 2496 2497 
    -- members (1) 
      -- 	branch_block_stmt_2042/merge_stmt_3907_PhiAck/$entry
      -- 
    cp_elements(2495) <= cp_elements(2494);
    -- CP-element group 2496 transition  input  bypass 
    -- predecessors 2495 
    -- successors 2498 
    -- members (1) 
      -- 	branch_block_stmt_2042/merge_stmt_3907_PhiAck/phi_stmt_3908_ack
      -- 
    phi_stmt_3908_ack_20178_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_3908_ack_0, ack => cp_elements(2496)); -- 
    -- CP-element group 2497 transition  input  bypass 
    -- predecessors 2495 
    -- successors 2498 
    -- members (1) 
      -- 	branch_block_stmt_2042/merge_stmt_3907_PhiAck/phi_stmt_3915_ack
      -- 
    phi_stmt_3915_ack_20179_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_3915_ack_0, ack => cp_elements(2497)); -- 
    -- CP-element group 2498 join  transition  bypass 
    -- predecessors 2496 2497 
    -- successors 75 
    -- members (1) 
      -- 	branch_block_stmt_2042/merge_stmt_3907_PhiAck/$exit
      -- 
    cp_element_group_2498: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_2498"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(2496) & cp_elements(2497);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(2498), clk => clk, reset => reset); --
    end block;
    -- CP-element group 2499 fork  transition  bypass 
    -- predecessors 1222 
    -- successors 2500 2506 
    -- members (1) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xi_udiv32x_xexitx_xx_xcritedge_crit_edgex_xi_PhiReq/$entry
      -- 
    cp_elements(2499) <= cp_elements(1222);
    -- CP-element group 2500 fork  transition  bypass 
    -- predecessors 2499 
    -- successors 2501 2503 
    -- members (4) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xi_udiv32x_xexitx_xx_xcritedge_crit_edgex_xi_PhiReq/phi_stmt_3966/$entry
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xi_udiv32x_xexitx_xx_xcritedge_crit_edgex_xi_PhiReq/phi_stmt_3966/phi_stmt_3966_sources/$entry
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xi_udiv32x_xexitx_xx_xcritedge_crit_edgex_xi_PhiReq/phi_stmt_3966/phi_stmt_3966_sources/type_cast_3969/$entry
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xi_udiv32x_xexitx_xx_xcritedge_crit_edgex_xi_PhiReq/phi_stmt_3966/phi_stmt_3966_sources/type_cast_3969/SplitProtocol/$entry
      -- 
    cp_elements(2500) <= cp_elements(2499);
    -- CP-element group 2501 transition  output  bypass 
    -- predecessors 2500 
    -- successors 2502 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xi_udiv32x_xexitx_xx_xcritedge_crit_edgex_xi_PhiReq/phi_stmt_3966/phi_stmt_3966_sources/type_cast_3969/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xi_udiv32x_xexitx_xx_xcritedge_crit_edgex_xi_PhiReq/phi_stmt_3966/phi_stmt_3966_sources/type_cast_3969/SplitProtocol/Sample/rr
      -- 
    cp_elements(2501) <= cp_elements(2500);
    rr_20202_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2501), ack => type_cast_3969_inst_req_0); -- 
    -- CP-element group 2502 transition  input  bypass 
    -- predecessors 2501 
    -- successors 2505 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xi_udiv32x_xexitx_xx_xcritedge_crit_edgex_xi_PhiReq/phi_stmt_3966/phi_stmt_3966_sources/type_cast_3969/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xi_udiv32x_xexitx_xx_xcritedge_crit_edgex_xi_PhiReq/phi_stmt_3966/phi_stmt_3966_sources/type_cast_3969/SplitProtocol/Sample/ra
      -- 
    ra_20203_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3969_inst_ack_0, ack => cp_elements(2502)); -- 
    -- CP-element group 2503 transition  output  bypass 
    -- predecessors 2500 
    -- successors 2504 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xi_udiv32x_xexitx_xx_xcritedge_crit_edgex_xi_PhiReq/phi_stmt_3966/phi_stmt_3966_sources/type_cast_3969/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xi_udiv32x_xexitx_xx_xcritedge_crit_edgex_xi_PhiReq/phi_stmt_3966/phi_stmt_3966_sources/type_cast_3969/SplitProtocol/Update/cr
      -- 
    cp_elements(2503) <= cp_elements(2500);
    cr_20207_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2503), ack => type_cast_3969_inst_req_1); -- 
    -- CP-element group 2504 transition  input  bypass 
    -- predecessors 2503 
    -- successors 2505 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xi_udiv32x_xexitx_xx_xcritedge_crit_edgex_xi_PhiReq/phi_stmt_3966/phi_stmt_3966_sources/type_cast_3969/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xi_udiv32x_xexitx_xx_xcritedge_crit_edgex_xi_PhiReq/phi_stmt_3966/phi_stmt_3966_sources/type_cast_3969/SplitProtocol/Update/ca
      -- 
    ca_20208_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3969_inst_ack_1, ack => cp_elements(2504)); -- 
    -- CP-element group 2505 join  transition  output  bypass 
    -- predecessors 2502 2504 
    -- successors 2512 
    -- members (5) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xi_udiv32x_xexitx_xx_xcritedge_crit_edgex_xi_PhiReq/phi_stmt_3966/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xi_udiv32x_xexitx_xx_xcritedge_crit_edgex_xi_PhiReq/phi_stmt_3966/phi_stmt_3966_sources/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xi_udiv32x_xexitx_xx_xcritedge_crit_edgex_xi_PhiReq/phi_stmt_3966/phi_stmt_3966_sources/type_cast_3969/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xi_udiv32x_xexitx_xx_xcritedge_crit_edgex_xi_PhiReq/phi_stmt_3966/phi_stmt_3966_sources/type_cast_3969/SplitProtocol/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xi_udiv32x_xexitx_xx_xcritedge_crit_edgex_xi_PhiReq/phi_stmt_3966/phi_stmt_3966_req
      -- 
    cp_element_group_2505: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_2505"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(2502) & cp_elements(2504);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(2505), clk => clk, reset => reset); --
    end block;
    phi_stmt_3966_req_20209_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2505), ack => phi_stmt_3966_req_0); -- 
    -- CP-element group 2506 fork  transition  bypass 
    -- predecessors 2499 
    -- successors 2507 2509 
    -- members (4) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xi_udiv32x_xexitx_xx_xcritedge_crit_edgex_xi_PhiReq/phi_stmt_3970/$entry
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xi_udiv32x_xexitx_xx_xcritedge_crit_edgex_xi_PhiReq/phi_stmt_3970/phi_stmt_3970_sources/$entry
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xi_udiv32x_xexitx_xx_xcritedge_crit_edgex_xi_PhiReq/phi_stmt_3970/phi_stmt_3970_sources/type_cast_3973/$entry
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xi_udiv32x_xexitx_xx_xcritedge_crit_edgex_xi_PhiReq/phi_stmt_3970/phi_stmt_3970_sources/type_cast_3973/SplitProtocol/$entry
      -- 
    cp_elements(2506) <= cp_elements(2499);
    -- CP-element group 2507 transition  output  bypass 
    -- predecessors 2506 
    -- successors 2508 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xi_udiv32x_xexitx_xx_xcritedge_crit_edgex_xi_PhiReq/phi_stmt_3970/phi_stmt_3970_sources/type_cast_3973/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xi_udiv32x_xexitx_xx_xcritedge_crit_edgex_xi_PhiReq/phi_stmt_3970/phi_stmt_3970_sources/type_cast_3973/SplitProtocol/Sample/rr
      -- 
    cp_elements(2507) <= cp_elements(2506);
    rr_20225_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2507), ack => type_cast_3973_inst_req_0); -- 
    -- CP-element group 2508 transition  input  bypass 
    -- predecessors 2507 
    -- successors 2511 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xi_udiv32x_xexitx_xx_xcritedge_crit_edgex_xi_PhiReq/phi_stmt_3970/phi_stmt_3970_sources/type_cast_3973/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xi_udiv32x_xexitx_xx_xcritedge_crit_edgex_xi_PhiReq/phi_stmt_3970/phi_stmt_3970_sources/type_cast_3973/SplitProtocol/Sample/ra
      -- 
    ra_20226_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3973_inst_ack_0, ack => cp_elements(2508)); -- 
    -- CP-element group 2509 transition  output  bypass 
    -- predecessors 2506 
    -- successors 2510 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xi_udiv32x_xexitx_xx_xcritedge_crit_edgex_xi_PhiReq/phi_stmt_3970/phi_stmt_3970_sources/type_cast_3973/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xi_udiv32x_xexitx_xx_xcritedge_crit_edgex_xi_PhiReq/phi_stmt_3970/phi_stmt_3970_sources/type_cast_3973/SplitProtocol/Update/cr
      -- 
    cp_elements(2509) <= cp_elements(2506);
    cr_20230_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2509), ack => type_cast_3973_inst_req_1); -- 
    -- CP-element group 2510 transition  input  bypass 
    -- predecessors 2509 
    -- successors 2511 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xi_udiv32x_xexitx_xx_xcritedge_crit_edgex_xi_PhiReq/phi_stmt_3970/phi_stmt_3970_sources/type_cast_3973/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xi_udiv32x_xexitx_xx_xcritedge_crit_edgex_xi_PhiReq/phi_stmt_3970/phi_stmt_3970_sources/type_cast_3973/SplitProtocol/Update/ca
      -- 
    ca_20231_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3973_inst_ack_1, ack => cp_elements(2510)); -- 
    -- CP-element group 2511 join  transition  output  bypass 
    -- predecessors 2508 2510 
    -- successors 2512 
    -- members (5) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xi_udiv32x_xexitx_xx_xcritedge_crit_edgex_xi_PhiReq/phi_stmt_3970/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xi_udiv32x_xexitx_xx_xcritedge_crit_edgex_xi_PhiReq/phi_stmt_3970/phi_stmt_3970_sources/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xi_udiv32x_xexitx_xx_xcritedge_crit_edgex_xi_PhiReq/phi_stmt_3970/phi_stmt_3970_sources/type_cast_3973/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xi_udiv32x_xexitx_xx_xcritedge_crit_edgex_xi_PhiReq/phi_stmt_3970/phi_stmt_3970_sources/type_cast_3973/SplitProtocol/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xi_udiv32x_xexitx_xx_xcritedge_crit_edgex_xi_PhiReq/phi_stmt_3970/phi_stmt_3970_req
      -- 
    cp_element_group_2511: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_2511"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(2508) & cp_elements(2510);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(2511), clk => clk, reset => reset); --
    end block;
    phi_stmt_3970_req_20232_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2511), ack => phi_stmt_3970_req_0); -- 
    -- CP-element group 2512 join  transition  bypass 
    -- predecessors 2505 2511 
    -- successors 2513 
    -- members (1) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xi_udiv32x_xexitx_xx_xcritedge_crit_edgex_xi_PhiReq/$exit
      -- 
    cp_element_group_2512: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_2512"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(2505) & cp_elements(2511);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(2512), clk => clk, reset => reset); --
    end block;
    -- CP-element group 2513 place  bypass 
    -- predecessors 2512 
    -- successors 2514 
    -- members (1) 
      -- 	branch_block_stmt_2042/merge_stmt_3965_PhiReqMerge
      -- 
    cp_elements(2513) <= cp_elements(2512);
    -- CP-element group 2514 fork  transition  bypass 
    -- predecessors 2513 
    -- successors 2515 2516 
    -- members (1) 
      -- 	branch_block_stmt_2042/merge_stmt_3965_PhiAck/$entry
      -- 
    cp_elements(2514) <= cp_elements(2513);
    -- CP-element group 2515 transition  input  bypass 
    -- predecessors 2514 
    -- successors 2517 
    -- members (1) 
      -- 	branch_block_stmt_2042/merge_stmt_3965_PhiAck/phi_stmt_3966_ack
      -- 
    phi_stmt_3966_ack_20237_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_3966_ack_0, ack => cp_elements(2515)); -- 
    -- CP-element group 2516 transition  input  bypass 
    -- predecessors 2514 
    -- successors 2517 
    -- members (1) 
      -- 	branch_block_stmt_2042/merge_stmt_3965_PhiAck/phi_stmt_3970_ack
      -- 
    phi_stmt_3970_ack_20238_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_3970_ack_0, ack => cp_elements(2516)); -- 
    -- CP-element group 2517 join  transition  bypass 
    -- predecessors 2515 2516 
    -- successors 77 
    -- members (1) 
      -- 	branch_block_stmt_2042/merge_stmt_3965_PhiAck/$exit
      -- 
    cp_element_group_2517: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_2517"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(2515) & cp_elements(2516);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(2517), clk => clk, reset => reset); --
    end block;
    -- CP-element group 2518 fork  transition  bypass 
    -- predecessors 1188 
    -- successors 2519 2531 
    -- members (1) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xpreheaderx_xi_xx_xcritedgex_xi_PhiReq/$entry
      -- 
    cp_elements(2518) <= cp_elements(1188);
    -- CP-element group 2519 fork  transition  bypass 
    -- predecessors 2518 
    -- successors 2520 2524 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xpreheaderx_xi_xx_xcritedgex_xi_PhiReq/phi_stmt_3988/$entry
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xpreheaderx_xi_xx_xcritedgex_xi_PhiReq/phi_stmt_3988/phi_stmt_3988_sources/$entry
      -- 
    cp_elements(2519) <= cp_elements(2518);
    -- CP-element group 2520 fork  transition  bypass 
    -- predecessors 2519 
    -- successors 2521 2522 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xpreheaderx_xi_xx_xcritedgex_xi_PhiReq/phi_stmt_3988/phi_stmt_3988_sources/type_cast_3991/$entry
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xpreheaderx_xi_xx_xcritedgex_xi_PhiReq/phi_stmt_3988/phi_stmt_3988_sources/type_cast_3991/SplitProtocol/$entry
      -- 
    cp_elements(2520) <= cp_elements(2519);
    -- CP-element group 2521 transition  bypass 
    -- predecessors 2520 
    -- successors 2523 
    -- members (4) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xpreheaderx_xi_xx_xcritedgex_xi_PhiReq/phi_stmt_3988/phi_stmt_3988_sources/type_cast_3991/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xpreheaderx_xi_xx_xcritedgex_xi_PhiReq/phi_stmt_3988/phi_stmt_3988_sources/type_cast_3991/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xpreheaderx_xi_xx_xcritedgex_xi_PhiReq/phi_stmt_3988/phi_stmt_3988_sources/type_cast_3991/SplitProtocol/Sample/rr
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xpreheaderx_xi_xx_xcritedgex_xi_PhiReq/phi_stmt_3988/phi_stmt_3988_sources/type_cast_3991/SplitProtocol/Sample/ra
      -- 
    cp_elements(2521) <= cp_elements(2520);
    -- CP-element group 2522 transition  bypass 
    -- predecessors 2520 
    -- successors 2523 
    -- members (4) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xpreheaderx_xi_xx_xcritedgex_xi_PhiReq/phi_stmt_3988/phi_stmt_3988_sources/type_cast_3991/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xpreheaderx_xi_xx_xcritedgex_xi_PhiReq/phi_stmt_3988/phi_stmt_3988_sources/type_cast_3991/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xpreheaderx_xi_xx_xcritedgex_xi_PhiReq/phi_stmt_3988/phi_stmt_3988_sources/type_cast_3991/SplitProtocol/Update/cr
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xpreheaderx_xi_xx_xcritedgex_xi_PhiReq/phi_stmt_3988/phi_stmt_3988_sources/type_cast_3991/SplitProtocol/Update/ca
      -- 
    cp_elements(2522) <= cp_elements(2520);
    -- CP-element group 2523 join  transition  bypass 
    -- predecessors 2521 2522 
    -- successors 2530 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xpreheaderx_xi_xx_xcritedgex_xi_PhiReq/phi_stmt_3988/phi_stmt_3988_sources/type_cast_3991/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xpreheaderx_xi_xx_xcritedgex_xi_PhiReq/phi_stmt_3988/phi_stmt_3988_sources/type_cast_3991/SplitProtocol/$exit
      -- 
    cp_element_group_2523: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_2523"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(2521) & cp_elements(2522);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(2523), clk => clk, reset => reset); --
    end block;
    -- CP-element group 2524 fork  transition  bypass 
    -- predecessors 2519 
    -- successors 2525 2527 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xpreheaderx_xi_xx_xcritedgex_xi_PhiReq/phi_stmt_3988/phi_stmt_3988_sources/type_cast_3993/$entry
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xpreheaderx_xi_xx_xcritedgex_xi_PhiReq/phi_stmt_3988/phi_stmt_3988_sources/type_cast_3993/SplitProtocol/$entry
      -- 
    cp_elements(2524) <= cp_elements(2519);
    -- CP-element group 2525 transition  output  bypass 
    -- predecessors 2524 
    -- successors 2526 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xpreheaderx_xi_xx_xcritedgex_xi_PhiReq/phi_stmt_3988/phi_stmt_3988_sources/type_cast_3993/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xpreheaderx_xi_xx_xcritedgex_xi_PhiReq/phi_stmt_3988/phi_stmt_3988_sources/type_cast_3993/SplitProtocol/Sample/rr
      -- 
    cp_elements(2525) <= cp_elements(2524);
    rr_20273_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2525), ack => type_cast_3993_inst_req_0); -- 
    -- CP-element group 2526 transition  input  bypass 
    -- predecessors 2525 
    -- successors 2529 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xpreheaderx_xi_xx_xcritedgex_xi_PhiReq/phi_stmt_3988/phi_stmt_3988_sources/type_cast_3993/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xpreheaderx_xi_xx_xcritedgex_xi_PhiReq/phi_stmt_3988/phi_stmt_3988_sources/type_cast_3993/SplitProtocol/Sample/ra
      -- 
    ra_20274_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3993_inst_ack_0, ack => cp_elements(2526)); -- 
    -- CP-element group 2527 transition  output  bypass 
    -- predecessors 2524 
    -- successors 2528 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xpreheaderx_xi_xx_xcritedgex_xi_PhiReq/phi_stmt_3988/phi_stmt_3988_sources/type_cast_3993/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xpreheaderx_xi_xx_xcritedgex_xi_PhiReq/phi_stmt_3988/phi_stmt_3988_sources/type_cast_3993/SplitProtocol/Update/cr
      -- 
    cp_elements(2527) <= cp_elements(2524);
    cr_20278_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2527), ack => type_cast_3993_inst_req_1); -- 
    -- CP-element group 2528 transition  input  bypass 
    -- predecessors 2527 
    -- successors 2529 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xpreheaderx_xi_xx_xcritedgex_xi_PhiReq/phi_stmt_3988/phi_stmt_3988_sources/type_cast_3993/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xpreheaderx_xi_xx_xcritedgex_xi_PhiReq/phi_stmt_3988/phi_stmt_3988_sources/type_cast_3993/SplitProtocol/Update/ca
      -- 
    ca_20279_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3993_inst_ack_1, ack => cp_elements(2528)); -- 
    -- CP-element group 2529 join  transition  bypass 
    -- predecessors 2526 2528 
    -- successors 2530 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xpreheaderx_xi_xx_xcritedgex_xi_PhiReq/phi_stmt_3988/phi_stmt_3988_sources/type_cast_3993/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xpreheaderx_xi_xx_xcritedgex_xi_PhiReq/phi_stmt_3988/phi_stmt_3988_sources/type_cast_3993/SplitProtocol/$exit
      -- 
    cp_element_group_2529: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_2529"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(2526) & cp_elements(2528);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(2529), clk => clk, reset => reset); --
    end block;
    -- CP-element group 2530 join  transition  output  bypass 
    -- predecessors 2523 2529 
    -- successors 2543 
    -- members (3) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xpreheaderx_xi_xx_xcritedgex_xi_PhiReq/phi_stmt_3988/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xpreheaderx_xi_xx_xcritedgex_xi_PhiReq/phi_stmt_3988/phi_stmt_3988_sources/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xpreheaderx_xi_xx_xcritedgex_xi_PhiReq/phi_stmt_3988/phi_stmt_3988_req
      -- 
    cp_element_group_2530: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_2530"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(2523) & cp_elements(2529);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(2530), clk => clk, reset => reset); --
    end block;
    phi_stmt_3988_req_20280_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2530), ack => phi_stmt_3988_req_1); -- 
    -- CP-element group 2531 fork  transition  bypass 
    -- predecessors 2518 
    -- successors 2532 2536 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xpreheaderx_xi_xx_xcritedgex_xi_PhiReq/phi_stmt_3994/$entry
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xpreheaderx_xi_xx_xcritedgex_xi_PhiReq/phi_stmt_3994/phi_stmt_3994_sources/$entry
      -- 
    cp_elements(2531) <= cp_elements(2518);
    -- CP-element group 2532 fork  transition  bypass 
    -- predecessors 2531 
    -- successors 2533 2534 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xpreheaderx_xi_xx_xcritedgex_xi_PhiReq/phi_stmt_3994/phi_stmt_3994_sources/type_cast_3997/$entry
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xpreheaderx_xi_xx_xcritedgex_xi_PhiReq/phi_stmt_3994/phi_stmt_3994_sources/type_cast_3997/SplitProtocol/$entry
      -- 
    cp_elements(2532) <= cp_elements(2531);
    -- CP-element group 2533 transition  bypass 
    -- predecessors 2532 
    -- successors 2535 
    -- members (4) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xpreheaderx_xi_xx_xcritedgex_xi_PhiReq/phi_stmt_3994/phi_stmt_3994_sources/type_cast_3997/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xpreheaderx_xi_xx_xcritedgex_xi_PhiReq/phi_stmt_3994/phi_stmt_3994_sources/type_cast_3997/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xpreheaderx_xi_xx_xcritedgex_xi_PhiReq/phi_stmt_3994/phi_stmt_3994_sources/type_cast_3997/SplitProtocol/Sample/rr
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xpreheaderx_xi_xx_xcritedgex_xi_PhiReq/phi_stmt_3994/phi_stmt_3994_sources/type_cast_3997/SplitProtocol/Sample/ra
      -- 
    cp_elements(2533) <= cp_elements(2532);
    -- CP-element group 2534 transition  bypass 
    -- predecessors 2532 
    -- successors 2535 
    -- members (4) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xpreheaderx_xi_xx_xcritedgex_xi_PhiReq/phi_stmt_3994/phi_stmt_3994_sources/type_cast_3997/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xpreheaderx_xi_xx_xcritedgex_xi_PhiReq/phi_stmt_3994/phi_stmt_3994_sources/type_cast_3997/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xpreheaderx_xi_xx_xcritedgex_xi_PhiReq/phi_stmt_3994/phi_stmt_3994_sources/type_cast_3997/SplitProtocol/Update/cr
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xpreheaderx_xi_xx_xcritedgex_xi_PhiReq/phi_stmt_3994/phi_stmt_3994_sources/type_cast_3997/SplitProtocol/Update/ca
      -- 
    cp_elements(2534) <= cp_elements(2532);
    -- CP-element group 2535 join  transition  bypass 
    -- predecessors 2533 2534 
    -- successors 2542 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xpreheaderx_xi_xx_xcritedgex_xi_PhiReq/phi_stmt_3994/phi_stmt_3994_sources/type_cast_3997/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xpreheaderx_xi_xx_xcritedgex_xi_PhiReq/phi_stmt_3994/phi_stmt_3994_sources/type_cast_3997/SplitProtocol/$exit
      -- 
    cp_element_group_2535: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_2535"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(2533) & cp_elements(2534);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(2535), clk => clk, reset => reset); --
    end block;
    -- CP-element group 2536 fork  transition  bypass 
    -- predecessors 2531 
    -- successors 2537 2539 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xpreheaderx_xi_xx_xcritedgex_xi_PhiReq/phi_stmt_3994/phi_stmt_3994_sources/type_cast_3999/$entry
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xpreheaderx_xi_xx_xcritedgex_xi_PhiReq/phi_stmt_3994/phi_stmt_3994_sources/type_cast_3999/SplitProtocol/$entry
      -- 
    cp_elements(2536) <= cp_elements(2531);
    -- CP-element group 2537 transition  output  bypass 
    -- predecessors 2536 
    -- successors 2538 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xpreheaderx_xi_xx_xcritedgex_xi_PhiReq/phi_stmt_3994/phi_stmt_3994_sources/type_cast_3999/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xpreheaderx_xi_xx_xcritedgex_xi_PhiReq/phi_stmt_3994/phi_stmt_3994_sources/type_cast_3999/SplitProtocol/Sample/rr
      -- 
    cp_elements(2537) <= cp_elements(2536);
    rr_20312_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2537), ack => type_cast_3999_inst_req_0); -- 
    -- CP-element group 2538 transition  input  bypass 
    -- predecessors 2537 
    -- successors 2541 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xpreheaderx_xi_xx_xcritedgex_xi_PhiReq/phi_stmt_3994/phi_stmt_3994_sources/type_cast_3999/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xpreheaderx_xi_xx_xcritedgex_xi_PhiReq/phi_stmt_3994/phi_stmt_3994_sources/type_cast_3999/SplitProtocol/Sample/ra
      -- 
    ra_20313_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3999_inst_ack_0, ack => cp_elements(2538)); -- 
    -- CP-element group 2539 transition  output  bypass 
    -- predecessors 2536 
    -- successors 2540 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xpreheaderx_xi_xx_xcritedgex_xi_PhiReq/phi_stmt_3994/phi_stmt_3994_sources/type_cast_3999/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xpreheaderx_xi_xx_xcritedgex_xi_PhiReq/phi_stmt_3994/phi_stmt_3994_sources/type_cast_3999/SplitProtocol/Update/cr
      -- 
    cp_elements(2539) <= cp_elements(2536);
    cr_20317_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2539), ack => type_cast_3999_inst_req_1); -- 
    -- CP-element group 2540 transition  input  bypass 
    -- predecessors 2539 
    -- successors 2541 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xpreheaderx_xi_xx_xcritedgex_xi_PhiReq/phi_stmt_3994/phi_stmt_3994_sources/type_cast_3999/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xpreheaderx_xi_xx_xcritedgex_xi_PhiReq/phi_stmt_3994/phi_stmt_3994_sources/type_cast_3999/SplitProtocol/Update/ca
      -- 
    ca_20318_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3999_inst_ack_1, ack => cp_elements(2540)); -- 
    -- CP-element group 2541 join  transition  bypass 
    -- predecessors 2538 2540 
    -- successors 2542 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xpreheaderx_xi_xx_xcritedgex_xi_PhiReq/phi_stmt_3994/phi_stmt_3994_sources/type_cast_3999/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xpreheaderx_xi_xx_xcritedgex_xi_PhiReq/phi_stmt_3994/phi_stmt_3994_sources/type_cast_3999/SplitProtocol/$exit
      -- 
    cp_element_group_2541: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_2541"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(2538) & cp_elements(2540);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(2541), clk => clk, reset => reset); --
    end block;
    -- CP-element group 2542 join  transition  output  bypass 
    -- predecessors 2535 2541 
    -- successors 2543 
    -- members (3) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xpreheaderx_xi_xx_xcritedgex_xi_PhiReq/phi_stmt_3994/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xpreheaderx_xi_xx_xcritedgex_xi_PhiReq/phi_stmt_3994/phi_stmt_3994_sources/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xpreheaderx_xi_xx_xcritedgex_xi_PhiReq/phi_stmt_3994/phi_stmt_3994_req
      -- 
    cp_element_group_2542: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_2542"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(2535) & cp_elements(2541);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(2542), clk => clk, reset => reset); --
    end block;
    phi_stmt_3994_req_20319_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2542), ack => phi_stmt_3994_req_1); -- 
    -- CP-element group 2543 join  transition  bypass 
    -- predecessors 2530 2542 
    -- successors 2570 
    -- members (1) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xpreheaderx_xi_xx_xcritedgex_xi_PhiReq/$exit
      -- 
    cp_element_group_2543: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_2543"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(2530) & cp_elements(2542);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(2543), clk => clk, reset => reset); --
    end block;
    -- CP-element group 2544 fork  transition  bypass 
    -- predecessors 1232 
    -- successors 2545 2557 
    -- members (1) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xx_xcritedge_crit_edgex_xi_xx_xcritedgex_xi_PhiReq/$entry
      -- 
    cp_elements(2544) <= cp_elements(1232);
    -- CP-element group 2545 fork  transition  bypass 
    -- predecessors 2544 
    -- successors 2546 2552 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xx_xcritedge_crit_edgex_xi_xx_xcritedgex_xi_PhiReq/phi_stmt_3988/$entry
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xx_xcritedge_crit_edgex_xi_xx_xcritedgex_xi_PhiReq/phi_stmt_3988/phi_stmt_3988_sources/$entry
      -- 
    cp_elements(2545) <= cp_elements(2544);
    -- CP-element group 2546 fork  transition  bypass 
    -- predecessors 2545 
    -- successors 2547 2549 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xx_xcritedge_crit_edgex_xi_xx_xcritedgex_xi_PhiReq/phi_stmt_3988/phi_stmt_3988_sources/type_cast_3991/$entry
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xx_xcritedge_crit_edgex_xi_xx_xcritedgex_xi_PhiReq/phi_stmt_3988/phi_stmt_3988_sources/type_cast_3991/SplitProtocol/$entry
      -- 
    cp_elements(2546) <= cp_elements(2545);
    -- CP-element group 2547 transition  output  bypass 
    -- predecessors 2546 
    -- successors 2548 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xx_xcritedge_crit_edgex_xi_xx_xcritedgex_xi_PhiReq/phi_stmt_3988/phi_stmt_3988_sources/type_cast_3991/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xx_xcritedge_crit_edgex_xi_xx_xcritedgex_xi_PhiReq/phi_stmt_3988/phi_stmt_3988_sources/type_cast_3991/SplitProtocol/Sample/rr
      -- 
    cp_elements(2547) <= cp_elements(2546);
    rr_20338_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2547), ack => type_cast_3991_inst_req_0); -- 
    -- CP-element group 2548 transition  input  bypass 
    -- predecessors 2547 
    -- successors 2551 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xx_xcritedge_crit_edgex_xi_xx_xcritedgex_xi_PhiReq/phi_stmt_3988/phi_stmt_3988_sources/type_cast_3991/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xx_xcritedge_crit_edgex_xi_xx_xcritedgex_xi_PhiReq/phi_stmt_3988/phi_stmt_3988_sources/type_cast_3991/SplitProtocol/Sample/ra
      -- 
    ra_20339_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3991_inst_ack_0, ack => cp_elements(2548)); -- 
    -- CP-element group 2549 transition  output  bypass 
    -- predecessors 2546 
    -- successors 2550 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xx_xcritedge_crit_edgex_xi_xx_xcritedgex_xi_PhiReq/phi_stmt_3988/phi_stmt_3988_sources/type_cast_3991/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xx_xcritedge_crit_edgex_xi_xx_xcritedgex_xi_PhiReq/phi_stmt_3988/phi_stmt_3988_sources/type_cast_3991/SplitProtocol/Update/cr
      -- 
    cp_elements(2549) <= cp_elements(2546);
    cr_20343_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2549), ack => type_cast_3991_inst_req_1); -- 
    -- CP-element group 2550 transition  input  bypass 
    -- predecessors 2549 
    -- successors 2551 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xx_xcritedge_crit_edgex_xi_xx_xcritedgex_xi_PhiReq/phi_stmt_3988/phi_stmt_3988_sources/type_cast_3991/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xx_xcritedge_crit_edgex_xi_xx_xcritedgex_xi_PhiReq/phi_stmt_3988/phi_stmt_3988_sources/type_cast_3991/SplitProtocol/Update/ca
      -- 
    ca_20344_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3991_inst_ack_1, ack => cp_elements(2550)); -- 
    -- CP-element group 2551 join  transition  bypass 
    -- predecessors 2548 2550 
    -- successors 2556 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xx_xcritedge_crit_edgex_xi_xx_xcritedgex_xi_PhiReq/phi_stmt_3988/phi_stmt_3988_sources/type_cast_3991/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xx_xcritedge_crit_edgex_xi_xx_xcritedgex_xi_PhiReq/phi_stmt_3988/phi_stmt_3988_sources/type_cast_3991/SplitProtocol/$exit
      -- 
    cp_element_group_2551: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_2551"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(2548) & cp_elements(2550);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(2551), clk => clk, reset => reset); --
    end block;
    -- CP-element group 2552 fork  transition  bypass 
    -- predecessors 2545 
    -- successors 2553 2554 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xx_xcritedge_crit_edgex_xi_xx_xcritedgex_xi_PhiReq/phi_stmt_3988/phi_stmt_3988_sources/type_cast_3993/$entry
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xx_xcritedge_crit_edgex_xi_xx_xcritedgex_xi_PhiReq/phi_stmt_3988/phi_stmt_3988_sources/type_cast_3993/SplitProtocol/$entry
      -- 
    cp_elements(2552) <= cp_elements(2545);
    -- CP-element group 2553 transition  bypass 
    -- predecessors 2552 
    -- successors 2555 
    -- members (4) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xx_xcritedge_crit_edgex_xi_xx_xcritedgex_xi_PhiReq/phi_stmt_3988/phi_stmt_3988_sources/type_cast_3993/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xx_xcritedge_crit_edgex_xi_xx_xcritedgex_xi_PhiReq/phi_stmt_3988/phi_stmt_3988_sources/type_cast_3993/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xx_xcritedge_crit_edgex_xi_xx_xcritedgex_xi_PhiReq/phi_stmt_3988/phi_stmt_3988_sources/type_cast_3993/SplitProtocol/Sample/rr
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xx_xcritedge_crit_edgex_xi_xx_xcritedgex_xi_PhiReq/phi_stmt_3988/phi_stmt_3988_sources/type_cast_3993/SplitProtocol/Sample/ra
      -- 
    cp_elements(2553) <= cp_elements(2552);
    -- CP-element group 2554 transition  bypass 
    -- predecessors 2552 
    -- successors 2555 
    -- members (4) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xx_xcritedge_crit_edgex_xi_xx_xcritedgex_xi_PhiReq/phi_stmt_3988/phi_stmt_3988_sources/type_cast_3993/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xx_xcritedge_crit_edgex_xi_xx_xcritedgex_xi_PhiReq/phi_stmt_3988/phi_stmt_3988_sources/type_cast_3993/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xx_xcritedge_crit_edgex_xi_xx_xcritedgex_xi_PhiReq/phi_stmt_3988/phi_stmt_3988_sources/type_cast_3993/SplitProtocol/Update/cr
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xx_xcritedge_crit_edgex_xi_xx_xcritedgex_xi_PhiReq/phi_stmt_3988/phi_stmt_3988_sources/type_cast_3993/SplitProtocol/Update/ca
      -- 
    cp_elements(2554) <= cp_elements(2552);
    -- CP-element group 2555 join  transition  bypass 
    -- predecessors 2553 2554 
    -- successors 2556 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xx_xcritedge_crit_edgex_xi_xx_xcritedgex_xi_PhiReq/phi_stmt_3988/phi_stmt_3988_sources/type_cast_3993/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xx_xcritedge_crit_edgex_xi_xx_xcritedgex_xi_PhiReq/phi_stmt_3988/phi_stmt_3988_sources/type_cast_3993/SplitProtocol/$exit
      -- 
    cp_element_group_2555: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_2555"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(2553) & cp_elements(2554);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(2555), clk => clk, reset => reset); --
    end block;
    -- CP-element group 2556 join  transition  output  bypass 
    -- predecessors 2551 2555 
    -- successors 2569 
    -- members (3) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xx_xcritedge_crit_edgex_xi_xx_xcritedgex_xi_PhiReq/phi_stmt_3988/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xx_xcritedge_crit_edgex_xi_xx_xcritedgex_xi_PhiReq/phi_stmt_3988/phi_stmt_3988_sources/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xx_xcritedge_crit_edgex_xi_xx_xcritedgex_xi_PhiReq/phi_stmt_3988/phi_stmt_3988_req
      -- 
    cp_element_group_2556: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_2556"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(2551) & cp_elements(2555);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(2556), clk => clk, reset => reset); --
    end block;
    phi_stmt_3988_req_20361_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2556), ack => phi_stmt_3988_req_0); -- 
    -- CP-element group 2557 fork  transition  bypass 
    -- predecessors 2544 
    -- successors 2558 2564 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xx_xcritedge_crit_edgex_xi_xx_xcritedgex_xi_PhiReq/phi_stmt_3994/$entry
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xx_xcritedge_crit_edgex_xi_xx_xcritedgex_xi_PhiReq/phi_stmt_3994/phi_stmt_3994_sources/$entry
      -- 
    cp_elements(2557) <= cp_elements(2544);
    -- CP-element group 2558 fork  transition  bypass 
    -- predecessors 2557 
    -- successors 2559 2561 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xx_xcritedge_crit_edgex_xi_xx_xcritedgex_xi_PhiReq/phi_stmt_3994/phi_stmt_3994_sources/type_cast_3997/$entry
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xx_xcritedge_crit_edgex_xi_xx_xcritedgex_xi_PhiReq/phi_stmt_3994/phi_stmt_3994_sources/type_cast_3997/SplitProtocol/$entry
      -- 
    cp_elements(2558) <= cp_elements(2557);
    -- CP-element group 2559 transition  output  bypass 
    -- predecessors 2558 
    -- successors 2560 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xx_xcritedge_crit_edgex_xi_xx_xcritedgex_xi_PhiReq/phi_stmt_3994/phi_stmt_3994_sources/type_cast_3997/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xx_xcritedge_crit_edgex_xi_xx_xcritedgex_xi_PhiReq/phi_stmt_3994/phi_stmt_3994_sources/type_cast_3997/SplitProtocol/Sample/rr
      -- 
    cp_elements(2559) <= cp_elements(2558);
    rr_20377_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2559), ack => type_cast_3997_inst_req_0); -- 
    -- CP-element group 2560 transition  input  bypass 
    -- predecessors 2559 
    -- successors 2563 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xx_xcritedge_crit_edgex_xi_xx_xcritedgex_xi_PhiReq/phi_stmt_3994/phi_stmt_3994_sources/type_cast_3997/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xx_xcritedge_crit_edgex_xi_xx_xcritedgex_xi_PhiReq/phi_stmt_3994/phi_stmt_3994_sources/type_cast_3997/SplitProtocol/Sample/ra
      -- 
    ra_20378_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3997_inst_ack_0, ack => cp_elements(2560)); -- 
    -- CP-element group 2561 transition  output  bypass 
    -- predecessors 2558 
    -- successors 2562 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xx_xcritedge_crit_edgex_xi_xx_xcritedgex_xi_PhiReq/phi_stmt_3994/phi_stmt_3994_sources/type_cast_3997/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xx_xcritedge_crit_edgex_xi_xx_xcritedgex_xi_PhiReq/phi_stmt_3994/phi_stmt_3994_sources/type_cast_3997/SplitProtocol/Update/cr
      -- 
    cp_elements(2561) <= cp_elements(2558);
    cr_20382_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2561), ack => type_cast_3997_inst_req_1); -- 
    -- CP-element group 2562 transition  input  bypass 
    -- predecessors 2561 
    -- successors 2563 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xx_xcritedge_crit_edgex_xi_xx_xcritedgex_xi_PhiReq/phi_stmt_3994/phi_stmt_3994_sources/type_cast_3997/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xx_xcritedge_crit_edgex_xi_xx_xcritedgex_xi_PhiReq/phi_stmt_3994/phi_stmt_3994_sources/type_cast_3997/SplitProtocol/Update/ca
      -- 
    ca_20383_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3997_inst_ack_1, ack => cp_elements(2562)); -- 
    -- CP-element group 2563 join  transition  bypass 
    -- predecessors 2560 2562 
    -- successors 2568 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xx_xcritedge_crit_edgex_xi_xx_xcritedgex_xi_PhiReq/phi_stmt_3994/phi_stmt_3994_sources/type_cast_3997/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xx_xcritedge_crit_edgex_xi_xx_xcritedgex_xi_PhiReq/phi_stmt_3994/phi_stmt_3994_sources/type_cast_3997/SplitProtocol/$exit
      -- 
    cp_element_group_2563: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_2563"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(2560) & cp_elements(2562);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(2563), clk => clk, reset => reset); --
    end block;
    -- CP-element group 2564 fork  transition  bypass 
    -- predecessors 2557 
    -- successors 2565 2566 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xx_xcritedge_crit_edgex_xi_xx_xcritedgex_xi_PhiReq/phi_stmt_3994/phi_stmt_3994_sources/type_cast_3999/$entry
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xx_xcritedge_crit_edgex_xi_xx_xcritedgex_xi_PhiReq/phi_stmt_3994/phi_stmt_3994_sources/type_cast_3999/SplitProtocol/$entry
      -- 
    cp_elements(2564) <= cp_elements(2557);
    -- CP-element group 2565 transition  bypass 
    -- predecessors 2564 
    -- successors 2567 
    -- members (4) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xx_xcritedge_crit_edgex_xi_xx_xcritedgex_xi_PhiReq/phi_stmt_3994/phi_stmt_3994_sources/type_cast_3999/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xx_xcritedge_crit_edgex_xi_xx_xcritedgex_xi_PhiReq/phi_stmt_3994/phi_stmt_3994_sources/type_cast_3999/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xx_xcritedge_crit_edgex_xi_xx_xcritedgex_xi_PhiReq/phi_stmt_3994/phi_stmt_3994_sources/type_cast_3999/SplitProtocol/Sample/rr
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xx_xcritedge_crit_edgex_xi_xx_xcritedgex_xi_PhiReq/phi_stmt_3994/phi_stmt_3994_sources/type_cast_3999/SplitProtocol/Sample/ra
      -- 
    cp_elements(2565) <= cp_elements(2564);
    -- CP-element group 2566 transition  bypass 
    -- predecessors 2564 
    -- successors 2567 
    -- members (4) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xx_xcritedge_crit_edgex_xi_xx_xcritedgex_xi_PhiReq/phi_stmt_3994/phi_stmt_3994_sources/type_cast_3999/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xx_xcritedge_crit_edgex_xi_xx_xcritedgex_xi_PhiReq/phi_stmt_3994/phi_stmt_3994_sources/type_cast_3999/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xx_xcritedge_crit_edgex_xi_xx_xcritedgex_xi_PhiReq/phi_stmt_3994/phi_stmt_3994_sources/type_cast_3999/SplitProtocol/Update/cr
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xx_xcritedge_crit_edgex_xi_xx_xcritedgex_xi_PhiReq/phi_stmt_3994/phi_stmt_3994_sources/type_cast_3999/SplitProtocol/Update/ca
      -- 
    cp_elements(2566) <= cp_elements(2564);
    -- CP-element group 2567 join  transition  bypass 
    -- predecessors 2565 2566 
    -- successors 2568 
    -- members (2) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xx_xcritedge_crit_edgex_xi_xx_xcritedgex_xi_PhiReq/phi_stmt_3994/phi_stmt_3994_sources/type_cast_3999/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xx_xcritedge_crit_edgex_xi_xx_xcritedgex_xi_PhiReq/phi_stmt_3994/phi_stmt_3994_sources/type_cast_3999/SplitProtocol/$exit
      -- 
    cp_element_group_2567: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_2567"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(2565) & cp_elements(2566);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(2567), clk => clk, reset => reset); --
    end block;
    -- CP-element group 2568 join  transition  output  bypass 
    -- predecessors 2563 2567 
    -- successors 2569 
    -- members (3) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xx_xcritedge_crit_edgex_xi_xx_xcritedgex_xi_PhiReq/phi_stmt_3994/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xx_xcritedge_crit_edgex_xi_xx_xcritedgex_xi_PhiReq/phi_stmt_3994/phi_stmt_3994_sources/$exit
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xx_xcritedge_crit_edgex_xi_xx_xcritedgex_xi_PhiReq/phi_stmt_3994/phi_stmt_3994_req
      -- 
    cp_element_group_2568: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_2568"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(2563) & cp_elements(2567);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(2568), clk => clk, reset => reset); --
    end block;
    phi_stmt_3994_req_20400_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2568), ack => phi_stmt_3994_req_0); -- 
    -- CP-element group 2569 join  transition  bypass 
    -- predecessors 2556 2568 
    -- successors 2570 
    -- members (1) 
      -- 	branch_block_stmt_2042/udiv32x_xexitx_xx_xcritedge_crit_edgex_xi_xx_xcritedgex_xi_PhiReq/$exit
      -- 
    cp_element_group_2569: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_2569"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(2556) & cp_elements(2568);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(2569), clk => clk, reset => reset); --
    end block;
    -- CP-element group 2570 merge  place  bypass 
    -- predecessors 2543 2569 
    -- successors 2571 
    -- members (1) 
      -- 	branch_block_stmt_2042/merge_stmt_3987_PhiReqMerge
      -- 
    cp_elements(2570) <= OrReduce(cp_elements(2543) & cp_elements(2569));
    -- CP-element group 2571 fork  transition  bypass 
    -- predecessors 2570 
    -- successors 2572 2573 
    -- members (1) 
      -- 	branch_block_stmt_2042/merge_stmt_3987_PhiAck/$entry
      -- 
    cp_elements(2571) <= cp_elements(2570);
    -- CP-element group 2572 transition  input  bypass 
    -- predecessors 2571 
    -- successors 2574 
    -- members (1) 
      -- 	branch_block_stmt_2042/merge_stmt_3987_PhiAck/phi_stmt_3988_ack
      -- 
    phi_stmt_3988_ack_20405_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_3988_ack_0, ack => cp_elements(2572)); -- 
    -- CP-element group 2573 transition  input  bypass 
    -- predecessors 2571 
    -- successors 2574 
    -- members (1) 
      -- 	branch_block_stmt_2042/merge_stmt_3987_PhiAck/phi_stmt_3994_ack
      -- 
    phi_stmt_3994_ack_20406_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_3994_ack_0, ack => cp_elements(2573)); -- 
    -- CP-element group 2574 join  transition  bypass 
    -- predecessors 2572 2573 
    -- successors 78 
    -- members (1) 
      -- 	branch_block_stmt_2042/merge_stmt_3987_PhiAck/$exit
      -- 
    cp_element_group_2574: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_2574"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(2572) & cp_elements(2573);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(2574), clk => clk, reset => reset); --
    end block;
    -- CP-element group 2575 transition  bypass 
    -- predecessors 1071 
    -- successors 2577 
    -- members (4) 
      -- 	branch_block_stmt_2042/bb_60_fdiv32x_xexit_PhiReq/phi_stmt_4035/phi_stmt_4035_sources/type_cast_4038/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_2042/bb_60_fdiv32x_xexit_PhiReq/phi_stmt_4035/phi_stmt_4035_sources/type_cast_4038/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_2042/bb_60_fdiv32x_xexit_PhiReq/phi_stmt_4035/phi_stmt_4035_sources/type_cast_4038/SplitProtocol/Sample/rr
      -- 	branch_block_stmt_2042/bb_60_fdiv32x_xexit_PhiReq/phi_stmt_4035/phi_stmt_4035_sources/type_cast_4038/SplitProtocol/Sample/ra
      -- 
    cp_elements(2575) <= cp_elements(1071);
    -- CP-element group 2576 transition  bypass 
    -- predecessors 1071 
    -- successors 2577 
    -- members (4) 
      -- 	branch_block_stmt_2042/bb_60_fdiv32x_xexit_PhiReq/phi_stmt_4035/phi_stmt_4035_sources/type_cast_4038/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_2042/bb_60_fdiv32x_xexit_PhiReq/phi_stmt_4035/phi_stmt_4035_sources/type_cast_4038/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_2042/bb_60_fdiv32x_xexit_PhiReq/phi_stmt_4035/phi_stmt_4035_sources/type_cast_4038/SplitProtocol/Update/cr
      -- 	branch_block_stmt_2042/bb_60_fdiv32x_xexit_PhiReq/phi_stmt_4035/phi_stmt_4035_sources/type_cast_4038/SplitProtocol/Update/ca
      -- 
    cp_elements(2576) <= cp_elements(1071);
    -- CP-element group 2577 join  transition  output  bypass 
    -- predecessors 2575 2576 
    -- successors 2583 
    -- members (6) 
      -- 	branch_block_stmt_2042/bb_60_fdiv32x_xexit_PhiReq/$exit
      -- 	branch_block_stmt_2042/bb_60_fdiv32x_xexit_PhiReq/phi_stmt_4035/$exit
      -- 	branch_block_stmt_2042/bb_60_fdiv32x_xexit_PhiReq/phi_stmt_4035/phi_stmt_4035_sources/$exit
      -- 	branch_block_stmt_2042/bb_60_fdiv32x_xexit_PhiReq/phi_stmt_4035/phi_stmt_4035_sources/type_cast_4038/$exit
      -- 	branch_block_stmt_2042/bb_60_fdiv32x_xexit_PhiReq/phi_stmt_4035/phi_stmt_4035_sources/type_cast_4038/SplitProtocol/$exit
      -- 	branch_block_stmt_2042/bb_60_fdiv32x_xexit_PhiReq/phi_stmt_4035/phi_stmt_4035_req
      -- 
    cp_element_group_2577: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_2577"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(2575) & cp_elements(2576);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(2577), clk => clk, reset => reset); --
    end block;
    phi_stmt_4035_req_20432_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2577), ack => phi_stmt_4035_req_1); -- 
    -- CP-element group 2578 transition  output  bypass 
    -- predecessors 1256 
    -- successors 2579 
    -- members (2) 
      -- 	branch_block_stmt_2042/xx_xcritedgex_xi_fdiv32x_xexit_PhiReq/phi_stmt_4035/phi_stmt_4035_sources/type_cast_4038/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_2042/xx_xcritedgex_xi_fdiv32x_xexit_PhiReq/phi_stmt_4035/phi_stmt_4035_sources/type_cast_4038/SplitProtocol/Sample/rr
      -- 
    cp_elements(2578) <= cp_elements(1256);
    rr_20451_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2578), ack => type_cast_4038_inst_req_0); -- 
    -- CP-element group 2579 transition  input  bypass 
    -- predecessors 2578 
    -- successors 2582 
    -- members (2) 
      -- 	branch_block_stmt_2042/xx_xcritedgex_xi_fdiv32x_xexit_PhiReq/phi_stmt_4035/phi_stmt_4035_sources/type_cast_4038/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_2042/xx_xcritedgex_xi_fdiv32x_xexit_PhiReq/phi_stmt_4035/phi_stmt_4035_sources/type_cast_4038/SplitProtocol/Sample/ra
      -- 
    ra_20452_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4038_inst_ack_0, ack => cp_elements(2579)); -- 
    -- CP-element group 2580 transition  output  bypass 
    -- predecessors 1256 
    -- successors 2581 
    -- members (2) 
      -- 	branch_block_stmt_2042/xx_xcritedgex_xi_fdiv32x_xexit_PhiReq/phi_stmt_4035/phi_stmt_4035_sources/type_cast_4038/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_2042/xx_xcritedgex_xi_fdiv32x_xexit_PhiReq/phi_stmt_4035/phi_stmt_4035_sources/type_cast_4038/SplitProtocol/Update/cr
      -- 
    cp_elements(2580) <= cp_elements(1256);
    cr_20456_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2580), ack => type_cast_4038_inst_req_1); -- 
    -- CP-element group 2581 transition  input  bypass 
    -- predecessors 2580 
    -- successors 2582 
    -- members (2) 
      -- 	branch_block_stmt_2042/xx_xcritedgex_xi_fdiv32x_xexit_PhiReq/phi_stmt_4035/phi_stmt_4035_sources/type_cast_4038/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_2042/xx_xcritedgex_xi_fdiv32x_xexit_PhiReq/phi_stmt_4035/phi_stmt_4035_sources/type_cast_4038/SplitProtocol/Update/ca
      -- 
    ca_20457_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4038_inst_ack_1, ack => cp_elements(2581)); -- 
    -- CP-element group 2582 join  transition  output  bypass 
    -- predecessors 2579 2581 
    -- successors 2583 
    -- members (6) 
      -- 	branch_block_stmt_2042/xx_xcritedgex_xi_fdiv32x_xexit_PhiReq/$exit
      -- 	branch_block_stmt_2042/xx_xcritedgex_xi_fdiv32x_xexit_PhiReq/phi_stmt_4035/$exit
      -- 	branch_block_stmt_2042/xx_xcritedgex_xi_fdiv32x_xexit_PhiReq/phi_stmt_4035/phi_stmt_4035_sources/$exit
      -- 	branch_block_stmt_2042/xx_xcritedgex_xi_fdiv32x_xexit_PhiReq/phi_stmt_4035/phi_stmt_4035_sources/type_cast_4038/$exit
      -- 	branch_block_stmt_2042/xx_xcritedgex_xi_fdiv32x_xexit_PhiReq/phi_stmt_4035/phi_stmt_4035_sources/type_cast_4038/SplitProtocol/$exit
      -- 	branch_block_stmt_2042/xx_xcritedgex_xi_fdiv32x_xexit_PhiReq/phi_stmt_4035/phi_stmt_4035_req
      -- 
    cp_element_group_2582: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_2582"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(2579) & cp_elements(2581);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(2582), clk => clk, reset => reset); --
    end block;
    phi_stmt_4035_req_20458_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2582), ack => phi_stmt_4035_req_0); -- 
    -- CP-element group 2583 merge  place  bypass 
    -- predecessors 2577 2582 
    -- successors 2584 
    -- members (1) 
      -- 	branch_block_stmt_2042/merge_stmt_4034_PhiReqMerge
      -- 
    cp_elements(2583) <= OrReduce(cp_elements(2577) & cp_elements(2582));
    -- CP-element group 2584 transition  bypass 
    -- predecessors 2583 
    -- successors 2585 
    -- members (1) 
      -- 	branch_block_stmt_2042/merge_stmt_4034_PhiAck/$entry
      -- 
    cp_elements(2584) <= cp_elements(2583);
    -- CP-element group 2585 transition  place  input  bypass 
    -- predecessors 2584 
    -- successors 1257 
    -- members (4) 
      -- 	branch_block_stmt_2042/merge_stmt_4034__exit__
      -- 	branch_block_stmt_2042/assign_stmt_4045__entry__
      -- 	branch_block_stmt_2042/merge_stmt_4034_PhiAck/$exit
      -- 	branch_block_stmt_2042/merge_stmt_4034_PhiAck/phi_stmt_4035_ack
      -- 
    phi_stmt_4035_ack_20463_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_4035_ack_0, ack => cp_elements(2585)); -- 
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal curr_quotientx_x02x_xix_xi_3764 : std_logic_vector(31 downto 0);
    signal curr_quotientx_x02x_xix_xix_xi35_2412 : std_logic_vector(31 downto 0);
    signal curr_quotientx_x02x_xix_xix_xi7_2853 : std_logic_vector(31 downto 0);
    signal curr_quotientx_x02x_xix_xix_xi_3299 : std_logic_vector(31 downto 0);
    signal curr_quotientx_x0x_xlcssax_xix_xi_3814 : std_logic_vector(31 downto 0);
    signal curr_quotientx_x0x_xlcssax_xix_xix_xi10_2902 : std_logic_vector(31 downto 0);
    signal curr_quotientx_x0x_xlcssax_xix_xix_xi38_2462 : std_logic_vector(31 downto 0);
    signal curr_quotientx_x0x_xlcssax_xix_xix_xi_3348 : std_logic_vector(31 downto 0);
    signal expr_2802_wire_constant : std_logic_vector(31 downto 0);
    signal expr_2802_wire_constant_cmp : std_logic_vector(0 downto 0);
    signal expr_2805_wire_constant : std_logic_vector(31 downto 0);
    signal expr_2805_wire_constant_cmp : std_logic_vector(0 downto 0);
    signal expr_3248_wire_constant : std_logic_vector(31 downto 0);
    signal expr_3248_wire_constant_cmp : std_logic_vector(0 downto 0);
    signal expr_3251_wire_constant : std_logic_vector(31 downto 0);
    signal expr_3251_wire_constant_cmp : std_logic_vector(0 downto 0);
    signal expx_x0x_xlcssax_xi_3988 : std_logic_vector(31 downto 0);
    signal expx_x0x_xlcssax_xix_xi25_3075 : std_logic_vector(31 downto 0);
    signal expx_x0x_xlcssax_xix_xi49_2636 : std_logic_vector(31 downto 0);
    signal expx_x0x_xlcssax_xix_xi_3521 : std_logic_vector(31 downto 0);
    signal flux_refx_x0_2304 : std_logic_vector(31 downto 0);
    signal flux_rotor_prevx_x0_2045 : std_logic_vector(31 downto 0);
    signal iNsTr_100_3245 : std_logic_vector(31 downto 0);
    signal iNsTr_104_2961 : std_logic_vector(31 downto 0);
    signal iNsTr_105_2967 : std_logic_vector(0 downto 0);
    signal iNsTr_106_2975 : std_logic_vector(0 downto 0);
    signal iNsTr_109_2474 : std_logic_vector(31 downto 0);
    signal iNsTr_10_2089 : std_logic_vector(31 downto 0);
    signal iNsTr_110_2479 : std_logic_vector(31 downto 0);
    signal iNsTr_111_2485 : std_logic_vector(0 downto 0);
    signal iNsTr_113_3642 : std_logic_vector(31 downto 0);
    signal iNsTr_114_3647 : std_logic_vector(31 downto 0);
    signal iNsTr_115_3653 : std_logic_vector(0 downto 0);
    signal iNsTr_117_3616 : std_logic_vector(0 downto 0);
    signal iNsTr_11_2094 : std_logic_vector(31 downto 0);
    signal iNsTr_121_3407 : std_logic_vector(31 downto 0);
    signal iNsTr_122_3413 : std_logic_vector(0 downto 0);
    signal iNsTr_123_3421 : std_logic_vector(0 downto 0);
    signal iNsTr_125_2832 : std_logic_vector(31 downto 0);
    signal iNsTr_126_2837 : std_logic_vector(0 downto 0);
    signal iNsTr_129_3093 : std_logic_vector(31 downto 0);
    signal iNsTr_12_2100 : std_logic_vector(31 downto 0);
    signal iNsTr_130_3099 : std_logic_vector(31 downto 0);
    signal iNsTr_131_3105 : std_logic_vector(31 downto 0);
    signal iNsTr_132_3110 : std_logic_vector(31 downto 0);
    signal iNsTr_133_3115 : std_logic_vector(31 downto 0);
    signal iNsTr_135_2425 : std_logic_vector(31 downto 0);
    signal iNsTr_136_2431 : std_logic_vector(31 downto 0);
    signal iNsTr_137_2436 : std_logic_vector(0 downto 0);
    signal iNsTr_139_2503 : std_logic_vector(31 downto 0);
    signal iNsTr_13_2105 : std_logic_vector(63 downto 0);
    signal iNsTr_140_2509 : std_logic_vector(31 downto 0);
    signal iNsTr_141_2515 : std_logic_vector(31 downto 0);
    signal iNsTr_142_2521 : std_logic_vector(31 downto 0);
    signal iNsTr_143_2527 : std_logic_vector(31 downto 0);
    signal iNsTr_144_2533 : std_logic_vector(0 downto 0);
    signal iNsTr_145_2541 : std_logic_vector(0 downto 0);
    signal iNsTr_147_3707 : std_logic_vector(31 downto 0);
    signal iNsTr_148_3713 : std_logic_vector(31 downto 0);
    signal iNsTr_149_3719 : std_logic_vector(31 downto 0);
    signal iNsTr_14_2111 : std_logic_vector(0 downto 0);
    signal iNsTr_151_3666 : std_logic_vector(0 downto 0);
    signal iNsTr_154_3278 : std_logic_vector(31 downto 0);
    signal iNsTr_155_3283 : std_logic_vector(0 downto 0);
    signal iNsTr_158_3539 : std_logic_vector(31 downto 0);
    signal iNsTr_159_3545 : std_logic_vector(31 downto 0);
    signal iNsTr_160_3551 : std_logic_vector(31 downto 0);
    signal iNsTr_161_3556 : std_logic_vector(31 downto 0);
    signal iNsTr_162_3561 : std_logic_vector(31 downto 0);
    signal iNsTr_165_2914 : std_logic_vector(31 downto 0);
    signal iNsTr_166_2919 : std_logic_vector(31 downto 0);
    signal iNsTr_167_2924 : std_logic_vector(0 downto 0);
    signal iNsTr_169_2990 : std_logic_vector(31 downto 0);
    signal iNsTr_16_2150 : std_logic_vector(31 downto 0);
    signal iNsTr_170_3009 : std_logic_vector(31 downto 0);
    signal iNsTr_171_3015 : std_logic_vector(31 downto 0);
    signal iNsTr_172_3021 : std_logic_vector(0 downto 0);
    signal iNsTr_173_3029 : std_logic_vector(0 downto 0);
    signal iNsTr_177_2654 : std_logic_vector(31 downto 0);
    signal iNsTr_178_2660 : std_logic_vector(31 downto 0);
    signal iNsTr_179_2666 : std_logic_vector(31 downto 0);
    signal iNsTr_17_2155 : std_logic_vector(31 downto 0);
    signal iNsTr_180_2671 : std_logic_vector(31 downto 0);
    signal iNsTr_181_2676 : std_logic_vector(31 downto 0);
    signal iNsTr_183_3741 : std_logic_vector(31 downto 0);
    signal iNsTr_184_3747 : std_logic_vector(0 downto 0);
    signal iNsTr_186_3679 : std_logic_vector(0 downto 0);
    signal iNsTr_189_3360 : std_logic_vector(31 downto 0);
    signal iNsTr_18_2161 : std_logic_vector(0 downto 0);
    signal iNsTr_190_3365 : std_logic_vector(31 downto 0);
    signal iNsTr_191_3370 : std_logic_vector(0 downto 0);
    signal iNsTr_193_3436 : std_logic_vector(31 downto 0);
    signal iNsTr_194_3455 : std_logic_vector(31 downto 0);
    signal iNsTr_195_3461 : std_logic_vector(31 downto 0);
    signal iNsTr_196_3467 : std_logic_vector(0 downto 0);
    signal iNsTr_197_3475 : std_logic_vector(0 downto 0);
    signal iNsTr_199_2866 : std_logic_vector(31 downto 0);
    signal iNsTr_200_2872 : std_logic_vector(31 downto 0);
    signal iNsTr_201_2877 : std_logic_vector(0 downto 0);
    signal iNsTr_205_2556 : std_logic_vector(31 downto 0);
    signal iNsTr_206_2575 : std_logic_vector(31 downto 0);
    signal iNsTr_207_2581 : std_logic_vector(31 downto 0);
    signal iNsTr_208_2587 : std_logic_vector(0 downto 0);
    signal iNsTr_209_2595 : std_logic_vector(0 downto 0);
    signal iNsTr_20_2124 : std_logic_vector(0 downto 0);
    signal iNsTr_212_3826 : std_logic_vector(31 downto 0);
    signal iNsTr_213_3831 : std_logic_vector(31 downto 0);
    signal iNsTr_214_3837 : std_logic_vector(0 downto 0);
    signal iNsTr_216_4035 : std_logic_vector(31 downto 0);
    signal iNsTr_226_3312 : std_logic_vector(31 downto 0);
    signal iNsTr_227_3318 : std_logic_vector(31 downto 0);
    signal iNsTr_228_3323 : std_logic_vector(0 downto 0);
    signal iNsTr_22_2204 : std_logic_vector(63 downto 0);
    signal iNsTr_234_3777 : std_logic_vector(31 downto 0);
    signal iNsTr_235_3783 : std_logic_vector(31 downto 0);
    signal iNsTr_236_3788 : std_logic_vector(0 downto 0);
    signal iNsTr_238_3855 : std_logic_vector(31 downto 0);
    signal iNsTr_239_3861 : std_logic_vector(31 downto 0);
    signal iNsTr_23_2210 : std_logic_vector(0 downto 0);
    signal iNsTr_240_3867 : std_logic_vector(31 downto 0);
    signal iNsTr_241_3873 : std_logic_vector(31 downto 0);
    signal iNsTr_242_3879 : std_logic_vector(31 downto 0);
    signal iNsTr_243_3885 : std_logic_vector(0 downto 0);
    signal iNsTr_244_3893 : std_logic_vector(0 downto 0);
    signal iNsTr_249_4006 : std_logic_vector(31 downto 0);
    signal iNsTr_250_4012 : std_logic_vector(31 downto 0);
    signal iNsTr_251_4018 : std_logic_vector(31 downto 0);
    signal iNsTr_252_4023 : std_logic_vector(31 downto 0);
    signal iNsTr_253_4028 : std_logic_vector(31 downto 0);
    signal iNsTr_255_3908 : std_logic_vector(31 downto 0);
    signal iNsTr_256_3927 : std_logic_vector(31 downto 0);
    signal iNsTr_257_3933 : std_logic_vector(31 downto 0);
    signal iNsTr_258_3939 : std_logic_vector(0 downto 0);
    signal iNsTr_259_3947 : std_logic_vector(0 downto 0);
    signal iNsTr_25_2174 : std_logic_vector(0 downto 0);
    signal iNsTr_28_2223 : std_logic_vector(0 downto 0);
    signal iNsTr_2_2069 : std_logic_vector(31 downto 0);
    signal iNsTr_30_2321 : std_logic_vector(31 downto 0);
    signal iNsTr_31_2327 : std_logic_vector(31 downto 0);
    signal iNsTr_32_2332 : std_logic_vector(31 downto 0);
    signal iNsTr_33_2342 : std_logic_vector(0 downto 0);
    signal iNsTr_36_2256 : std_logic_vector(0 downto 0);
    signal iNsTr_38_2236 : std_logic_vector(31 downto 0);
    signal iNsTr_39_2242 : std_logic_vector(31 downto 0);
    signal iNsTr_40_2248 : std_logic_vector(31 downto 0);
    signal iNsTr_42_2683 : std_logic_vector(31 downto 0);
    signal iNsTr_43_2696 : std_logic_vector(31 downto 0);
    signal iNsTr_44_2702 : std_logic_vector(31 downto 0);
    signal iNsTr_45_2716 : std_logic_vector(0 downto 0);
    signal iNsTr_47_2355 : std_logic_vector(31 downto 0);
    signal iNsTr_48_2361 : std_logic_vector(31 downto 0);
    signal iNsTr_49_2367 : std_logic_vector(31 downto 0);
    signal iNsTr_4_2072 : std_logic_vector(31 downto 0);
    signal iNsTr_51_2289 : std_logic_vector(31 downto 0);
    signal iNsTr_52_2295 : std_logic_vector(31 downto 0);
    signal iNsTr_53_2301 : std_logic_vector(31 downto 0);
    signal iNsTr_55_2269 : std_logic_vector(31 downto 0);
    signal iNsTr_56_2275 : std_logic_vector(31 downto 0);
    signal iNsTr_57_2281 : std_logic_vector(31 downto 0);
    signal iNsTr_59_3122 : std_logic_vector(31 downto 0);
    signal iNsTr_60_3135 : std_logic_vector(0 downto 0);
    signal iNsTr_61_3149 : std_logic_vector(31 downto 0);
    signal iNsTr_62_3162 : std_logic_vector(0 downto 0);
    signal iNsTr_64_2729 : std_logic_vector(31 downto 0);
    signal iNsTr_65_2735 : std_logic_vector(31 downto 0);
    signal iNsTr_66_2741 : std_logic_vector(31 downto 0);
    signal iNsTr_67_2747 : std_logic_vector(31 downto 0);
    signal iNsTr_68_2753 : std_logic_vector(31 downto 0);
    signal iNsTr_69_2759 : std_logic_vector(31 downto 0);
    signal iNsTr_6_2075 : std_logic_vector(31 downto 0);
    signal iNsTr_70_2765 : std_logic_vector(31 downto 0);
    signal iNsTr_71_2771 : std_logic_vector(31 downto 0);
    signal iNsTr_72_2777 : std_logic_vector(31 downto 0);
    signal iNsTr_73_2783 : std_logic_vector(31 downto 0);
    signal iNsTr_74_2788 : std_logic_vector(31 downto 0);
    signal iNsTr_75_2794 : std_logic_vector(31 downto 0);
    signal iNsTr_76_2799 : std_logic_vector(31 downto 0);
    signal iNsTr_78_2389 : std_logic_vector(31 downto 0);
    signal iNsTr_79_2395 : std_logic_vector(0 downto 0);
    signal iNsTr_81_3568 : std_logic_vector(31 downto 0);
    signal iNsTr_82_3580 : std_logic_vector(31 downto 0);
    signal iNsTr_83_3586 : std_logic_vector(31 downto 0);
    signal iNsTr_84_3591 : std_logic_vector(31 downto 0);
    signal iNsTr_85_3597 : std_logic_vector(31 downto 0);
    signal iNsTr_86_3603 : std_logic_vector(0 downto 0);
    signal iNsTr_88_3175 : std_logic_vector(31 downto 0);
    signal iNsTr_89_3181 : std_logic_vector(31 downto 0);
    signal iNsTr_8_2078 : std_logic_vector(31 downto 0);
    signal iNsTr_90_3187 : std_logic_vector(31 downto 0);
    signal iNsTr_91_3193 : std_logic_vector(31 downto 0);
    signal iNsTr_92_3199 : std_logic_vector(31 downto 0);
    signal iNsTr_93_3205 : std_logic_vector(31 downto 0);
    signal iNsTr_94_3211 : std_logic_vector(31 downto 0);
    signal iNsTr_95_3217 : std_logic_vector(31 downto 0);
    signal iNsTr_96_3223 : std_logic_vector(31 downto 0);
    signal iNsTr_97_3229 : std_logic_vector(31 downto 0);
    signal iNsTr_98_3234 : std_logic_vector(31 downto 0);
    signal iNsTr_99_3240 : std_logic_vector(31 downto 0);
    signal iNsTr_9_2083 : std_logic_vector(31 downto 0);
    signal indvarx_xnextx_xi_3958 : std_logic_vector(31 downto 0);
    signal indvarx_xnextx_xix_xi19_3040 : std_logic_vector(31 downto 0);
    signal indvarx_xnextx_xix_xi44_2606 : std_logic_vector(31 downto 0);
    signal indvarx_xnextx_xix_xi_3486 : std_logic_vector(31 downto 0);
    signal int_flux_errx_x0_2052 : std_logic_vector(31 downto 0);
    signal int_flux_errx_x1_3626 : std_logic_vector(31 downto 0);
    signal int_speed_errx_x0_2059 : std_logic_vector(31 downto 0);
    signal int_speed_errx_x1_2134 : std_logic_vector(31 downto 0);
    signal orx_xcond11x_xi_3898 : std_logic_vector(0 downto 0);
    signal orx_xcond11x_xix_xi15_2980 : std_logic_vector(0 downto 0);
    signal orx_xcond11x_xix_xi40_2546 : std_logic_vector(0 downto 0);
    signal orx_xcond11x_xix_xi_3426 : std_logic_vector(0 downto 0);
    signal orx_xcondx_xi_3952 : std_logic_vector(0 downto 0);
    signal orx_xcondx_xix_xi18_3034 : std_logic_vector(0 downto 0);
    signal orx_xcondx_xix_xi43_2600 : std_logic_vector(0 downto 0);
    signal orx_xcondx_xix_xi_3480 : std_logic_vector(0 downto 0);
    signal phitmp_2187 : std_logic_vector(31 downto 0);
    signal quotientx_x05x_xix_xi_3728 : std_logic_vector(31 downto 0);
    signal quotientx_x05x_xix_xix_xi32_2376 : std_logic_vector(31 downto 0);
    signal quotientx_x05x_xix_xix_xi4_2819 : std_logic_vector(31 downto 0);
    signal quotientx_x05x_xix_xix_xi_3265 : std_logic_vector(31 downto 0);
    signal shifted_divisorx_x03x_xix_xi_3757 : std_logic_vector(31 downto 0);
    signal shifted_divisorx_x03x_xix_xix_xi34_2405 : std_logic_vector(31 downto 0);
    signal shifted_divisorx_x03x_xix_xix_xi6_2847 : std_logic_vector(31 downto 0);
    signal shifted_divisorx_x03x_xix_xix_xi_3293 : std_logic_vector(31 downto 0);
    signal shifted_divisorx_x0x_xlcssax_xix_xi_3807 : std_logic_vector(31 downto 0);
    signal shifted_divisorx_x0x_xlcssax_xix_xix_xi37_2455 : std_logic_vector(31 downto 0);
    signal shifted_divisorx_x0x_xlcssax_xix_xix_xi9_2896 : std_logic_vector(31 downto 0);
    signal shifted_divisorx_x0x_xlcssax_xix_xix_xi_3342 : std_logic_vector(31 downto 0);
    signal tempx_x012x_xi_3915 : std_logic_vector(31 downto 0);
    signal tempx_x012x_xix_xi17_2997 : std_logic_vector(31 downto 0);
    signal tempx_x012x_xix_xi42_2563 : std_logic_vector(31 downto 0);
    signal tempx_x012x_xix_xi_3443 : std_logic_vector(31 downto 0);
    signal tempx_x0x_xlcssax_xi_3994 : std_logic_vector(31 downto 0);
    signal tempx_x0x_xlcssax_xix_xi26_3081 : std_logic_vector(31 downto 0);
    signal tempx_x0x_xlcssax_xix_xi50_2642 : std_logic_vector(31 downto 0);
    signal tempx_x0x_xlcssax_xix_xi_3527 : std_logic_vector(31 downto 0);
    signal tempx_x0x_xphx_xix_xi14_2949 : std_logic_vector(31 downto 0);
    signal tempx_x0x_xphx_xix_xi_3395 : std_logic_vector(31 downto 0);
    signal tmp10x_xi55_3701 : std_logic_vector(31 downto 0);
    signal tmp10x_xi55x_xin_3687 : std_logic_vector(31 downto 0);
    signal tmp10x_xix_xi1_2706 : std_logic_vector(31 downto 0);
    signal tmp10x_xix_xi30_2336 : std_logic_vector(31 downto 0);
    signal tmp10x_xix_xi_3145 : std_logic_vector(31 downto 0);
    signal tmp21x_xix_xi21_3062 : std_logic_vector(31 downto 0);
    signal tmp21x_xix_xi_3508 : std_logic_vector(31 downto 0);
    signal tmp25x_xi_3980 : std_logic_vector(31 downto 0);
    signal tmp25x_xix_xi22_3067 : std_logic_vector(31 downto 0);
    signal tmp25x_xix_xi46_2628 : std_logic_vector(31 downto 0);
    signal tmp25x_xix_xi_3513 : std_logic_vector(31 downto 0);
    signal tmp26x_xi_3985 : std_logic_vector(31 downto 0);
    signal tmp26x_xix_xi23_3072 : std_logic_vector(31 downto 0);
    signal tmp26x_xix_xi47_2633 : std_logic_vector(31 downto 0);
    signal tmp26x_xix_xi_3518 : std_logic_vector(31 downto 0);
    signal tmp3x_xi_4032 : std_logic_vector(31 downto 0);
    signal tmp3x_xix_xi27_3119 : std_logic_vector(31 downto 0);
    signal tmp3x_xix_xi51_2680 : std_logic_vector(31 downto 0);
    signal tmp3x_xix_xi_3565 : std_logic_vector(31 downto 0);
    signal tmp6x_xix_xi2_2710 : std_logic_vector(31 downto 0);
    signal tmp6x_xix_xi_3156 : std_logic_vector(31 downto 0);
    signal torque_refx_x0_2190 : std_logic_vector(31 downto 0);
    signal type_cast_2049_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2051_wire : std_logic_vector(31 downto 0);
    signal type_cast_2056_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2058_wire : std_logic_vector(31 downto 0);
    signal type_cast_2063_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2065_wire : std_logic_vector(31 downto 0);
    signal type_cast_2087_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2098_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2109_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2122_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2137_wire : std_logic_vector(31 downto 0);
    signal type_cast_2140_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2143_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2148_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2159_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2172_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2185_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2193_wire : std_logic_vector(31 downto 0);
    signal type_cast_2196_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2199_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2208_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2221_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2234_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2240_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2246_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2254_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2267_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2273_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2279_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2287_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2293_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2299_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2307_wire : std_logic_vector(31 downto 0);
    signal type_cast_2309_wire : std_logic_vector(31 downto 0);
    signal type_cast_2311_wire : std_logic_vector(31 downto 0);
    signal type_cast_2314_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2319_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2325_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2340_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2353_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2359_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2365_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2373_wire : std_logic_vector(31 downto 0);
    signal type_cast_2375_wire : std_logic_vector(31 downto 0);
    signal type_cast_2379_wire : std_logic_vector(31 downto 0);
    signal type_cast_2382_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2387_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2393_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2408_wire : std_logic_vector(31 downto 0);
    signal type_cast_2411_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2415_wire : std_logic_vector(31 downto 0);
    signal type_cast_2418_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2423_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2429_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2447_wire : std_logic_vector(31 downto 0);
    signal type_cast_2451_wire : std_logic_vector(31 downto 0);
    signal type_cast_2459_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2461_wire : std_logic_vector(31 downto 0);
    signal type_cast_2466_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2468_wire : std_logic_vector(31 downto 0);
    signal type_cast_2483_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2496_wire : std_logic_vector(31 downto 0);
    signal type_cast_2501_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2507_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2513_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2519_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2525_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2531_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2536_wire : std_logic_vector(31 downto 0);
    signal type_cast_2539_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2559_wire : std_logic_vector(31 downto 0);
    signal type_cast_2562_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2566_wire : std_logic_vector(31 downto 0);
    signal type_cast_2568_wire : std_logic_vector(31 downto 0);
    signal type_cast_2573_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2579_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2585_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2590_wire : std_logic_vector(31 downto 0);
    signal type_cast_2593_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2604_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2617_wire : std_logic_vector(31 downto 0);
    signal type_cast_2621_wire : std_logic_vector(31 downto 0);
    signal type_cast_2626_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2639_wire : std_logic_vector(31 downto 0);
    signal type_cast_2641_wire : std_logic_vector(31 downto 0);
    signal type_cast_2645_wire : std_logic_vector(31 downto 0);
    signal type_cast_2647_wire : std_logic_vector(31 downto 0);
    signal type_cast_2652_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2658_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2664_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2686_wire : std_logic_vector(31 downto 0);
    signal type_cast_2689_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2694_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2700_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2714_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2727_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2733_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2739_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2745_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2751_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2757_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2763_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2769_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2775_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2781_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2792_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2816_wire : std_logic_vector(31 downto 0);
    signal type_cast_2818_wire : std_logic_vector(31 downto 0);
    signal type_cast_2822_wire : std_logic_vector(31 downto 0);
    signal type_cast_2825_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2830_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2850_wire : std_logic_vector(31 downto 0);
    signal type_cast_2852_wire : std_logic_vector(31 downto 0);
    signal type_cast_2856_wire : std_logic_vector(31 downto 0);
    signal type_cast_2859_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2864_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2870_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2888_wire : std_logic_vector(31 downto 0);
    signal type_cast_2892_wire : std_logic_vector(31 downto 0);
    signal type_cast_2899_wire : std_logic_vector(31 downto 0);
    signal type_cast_2901_wire : std_logic_vector(31 downto 0);
    signal type_cast_2906_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2908_wire : std_logic_vector(31 downto 0);
    signal type_cast_2935_wire : std_logic_vector(31 downto 0);
    signal type_cast_2943_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2945_wire : std_logic_vector(31 downto 0);
    signal type_cast_2952_wire : std_logic_vector(31 downto 0);
    signal type_cast_2954_wire : std_logic_vector(31 downto 0);
    signal type_cast_2959_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2965_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2970_wire : std_logic_vector(31 downto 0);
    signal type_cast_2973_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2993_wire : std_logic_vector(31 downto 0);
    signal type_cast_2996_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3000_wire : std_logic_vector(31 downto 0);
    signal type_cast_3002_wire : std_logic_vector(31 downto 0);
    signal type_cast_3007_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3013_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3019_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3024_wire : std_logic_vector(31 downto 0);
    signal type_cast_3027_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3038_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3051_wire : std_logic_vector(31 downto 0);
    signal type_cast_3055_wire : std_logic_vector(31 downto 0);
    signal type_cast_3060_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3078_wire : std_logic_vector(31 downto 0);
    signal type_cast_3080_wire : std_logic_vector(31 downto 0);
    signal type_cast_3084_wire : std_logic_vector(31 downto 0);
    signal type_cast_3086_wire : std_logic_vector(31 downto 0);
    signal type_cast_3091_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3097_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3103_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3125_wire : std_logic_vector(31 downto 0);
    signal type_cast_3128_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3133_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3139_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3153_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3160_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3173_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3179_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3185_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3191_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3197_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3203_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3209_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3215_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3221_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3227_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3238_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3262_wire : std_logic_vector(31 downto 0);
    signal type_cast_3264_wire : std_logic_vector(31 downto 0);
    signal type_cast_3268_wire : std_logic_vector(31 downto 0);
    signal type_cast_3271_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3276_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3296_wire : std_logic_vector(31 downto 0);
    signal type_cast_3298_wire : std_logic_vector(31 downto 0);
    signal type_cast_3302_wire : std_logic_vector(31 downto 0);
    signal type_cast_3305_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3310_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3316_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3334_wire : std_logic_vector(31 downto 0);
    signal type_cast_3338_wire : std_logic_vector(31 downto 0);
    signal type_cast_3345_wire : std_logic_vector(31 downto 0);
    signal type_cast_3347_wire : std_logic_vector(31 downto 0);
    signal type_cast_3352_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3354_wire : std_logic_vector(31 downto 0);
    signal type_cast_3381_wire : std_logic_vector(31 downto 0);
    signal type_cast_3389_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3391_wire : std_logic_vector(31 downto 0);
    signal type_cast_3398_wire : std_logic_vector(31 downto 0);
    signal type_cast_3400_wire : std_logic_vector(31 downto 0);
    signal type_cast_3405_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3411_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3416_wire : std_logic_vector(31 downto 0);
    signal type_cast_3419_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3439_wire : std_logic_vector(31 downto 0);
    signal type_cast_3442_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3446_wire : std_logic_vector(31 downto 0);
    signal type_cast_3448_wire : std_logic_vector(31 downto 0);
    signal type_cast_3453_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3459_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3465_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3470_wire : std_logic_vector(31 downto 0);
    signal type_cast_3473_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3484_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3497_wire : std_logic_vector(31 downto 0);
    signal type_cast_3501_wire : std_logic_vector(31 downto 0);
    signal type_cast_3506_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3524_wire : std_logic_vector(31 downto 0);
    signal type_cast_3526_wire : std_logic_vector(31 downto 0);
    signal type_cast_3530_wire : std_logic_vector(31 downto 0);
    signal type_cast_3532_wire : std_logic_vector(31 downto 0);
    signal type_cast_3537_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3543_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3549_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3571_wire : std_logic_vector(31 downto 0);
    signal type_cast_3574_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3584_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3595_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3601_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3614_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3629_wire : std_logic_vector(31 downto 0);
    signal type_cast_3632_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3635_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3640_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3651_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3664_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3677_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3690_wire : std_logic_vector(31 downto 0);
    signal type_cast_3693_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3696_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3705_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3711_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3717_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3725_wire : std_logic_vector(31 downto 0);
    signal type_cast_3727_wire : std_logic_vector(31 downto 0);
    signal type_cast_3731_wire : std_logic_vector(31 downto 0);
    signal type_cast_3734_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3739_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3745_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3760_wire : std_logic_vector(31 downto 0);
    signal type_cast_3763_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3767_wire : std_logic_vector(31 downto 0);
    signal type_cast_3770_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3775_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3781_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3799_wire : std_logic_vector(31 downto 0);
    signal type_cast_3803_wire : std_logic_vector(31 downto 0);
    signal type_cast_3811_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3813_wire : std_logic_vector(31 downto 0);
    signal type_cast_3818_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3820_wire : std_logic_vector(31 downto 0);
    signal type_cast_3835_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3848_wire : std_logic_vector(31 downto 0);
    signal type_cast_3853_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3859_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3865_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3871_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3877_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3883_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3888_wire : std_logic_vector(31 downto 0);
    signal type_cast_3891_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3911_wire : std_logic_vector(31 downto 0);
    signal type_cast_3914_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3918_wire : std_logic_vector(31 downto 0);
    signal type_cast_3920_wire : std_logic_vector(31 downto 0);
    signal type_cast_3925_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3931_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3937_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3942_wire : std_logic_vector(31 downto 0);
    signal type_cast_3945_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3956_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3969_wire : std_logic_vector(31 downto 0);
    signal type_cast_3973_wire : std_logic_vector(31 downto 0);
    signal type_cast_3978_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3991_wire : std_logic_vector(31 downto 0);
    signal type_cast_3993_wire : std_logic_vector(31 downto 0);
    signal type_cast_3997_wire : std_logic_vector(31 downto 0);
    signal type_cast_3999_wire : std_logic_vector(31 downto 0);
    signal type_cast_4004_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_4010_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_4016_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_4038_wire : std_logic_vector(31 downto 0);
    signal type_cast_4041_wire_constant : std_logic_vector(31 downto 0);
    signal xx_x016x_xix_xi_3722 : std_logic_vector(31 downto 0);
    signal xx_x016x_xix_xix_xi31_2370 : std_logic_vector(31 downto 0);
    signal xx_x016x_xix_xix_xi3_2813 : std_logic_vector(31 downto 0);
    signal xx_x016x_xix_xix_xi_3259 : std_logic_vector(31 downto 0);
    signal xx_x0x_xix_xix_xi12_2939 : std_logic_vector(31 downto 0);
    signal xx_x0x_xix_xix_xi_3385 : std_logic_vector(31 downto 0);
    signal xx_xlcssa10_3052 : std_logic_vector(31 downto 0);
    signal xx_xlcssa11_3048 : std_logic_vector(31 downto 0);
    signal xx_xlcssa12_2889 : std_logic_vector(31 downto 0);
    signal xx_xlcssa13_2885 : std_logic_vector(31 downto 0);
    signal xx_xlcssa14_2932 : std_logic_vector(31 downto 0);
    signal xx_xlcssa15_2618 : std_logic_vector(31 downto 0);
    signal xx_xlcssa16_2614 : std_logic_vector(31 downto 0);
    signal xx_xlcssa17_2448 : std_logic_vector(31 downto 0);
    signal xx_xlcssa18_2444 : std_logic_vector(31 downto 0);
    signal xx_xlcssa19_2493 : std_logic_vector(31 downto 0);
    signal xx_xlcssa1_3966 : std_logic_vector(31 downto 0);
    signal xx_xlcssa2_3800 : std_logic_vector(31 downto 0);
    signal xx_xlcssa3_3796 : std_logic_vector(31 downto 0);
    signal xx_xlcssa4_3845 : std_logic_vector(31 downto 0);
    signal xx_xlcssa5_3498 : std_logic_vector(31 downto 0);
    signal xx_xlcssa6_3494 : std_logic_vector(31 downto 0);
    signal xx_xlcssa7_3335 : std_logic_vector(31 downto 0);
    signal xx_xlcssa8_3331 : std_logic_vector(31 downto 0);
    signal xx_xlcssa9_3378 : std_logic_vector(31 downto 0);
    signal xx_xlcssa_3970 : std_logic_vector(31 downto 0);
    signal xx_xop_3141 : std_logic_vector(31 downto 0);
    -- 
  begin -- 
    expr_2802_wire_constant <= "00000000000000000000000000000000";
    expr_2805_wire_constant <= "00000000000000000000000000000001";
    expr_3248_wire_constant <= "00000000000000000000000000000000";
    expr_3251_wire_constant <= "00000000000000000000000000000001";
    type_cast_2049_wire_constant <= "00000000000000000000000000000000";
    type_cast_2056_wire_constant <= "00000000000000000000000000000000";
    type_cast_2063_wire_constant <= "00000000000000000000000000000000";
    type_cast_2087_wire_constant <= "00111000010100011011011100010111";
    type_cast_2098_wire_constant <= "01000010010010000000000000000000";
    type_cast_2109_wire_constant <= "1100000000101110000000000000000000000000000000000000000000000000";
    type_cast_2122_wire_constant <= "0100000000101110000000000000000000000000000000000000000000000000";
    type_cast_2140_wire_constant <= "11000001011100000000000000000000";
    type_cast_2143_wire_constant <= "01000001011100000000000000000000";
    type_cast_2148_wire_constant <= "01000010001000000000000000000000";
    type_cast_2159_wire_constant <= "11000001111100000000000000000000";
    type_cast_2172_wire_constant <= "01000001111100000000000000000000";
    type_cast_2185_wire_constant <= "01000100110100100111000000000000";
    type_cast_2196_wire_constant <= "11000111010001010100100100000000";
    type_cast_2199_wire_constant <= "01000111010001010100100100000000";
    type_cast_2208_wire_constant <= "0100000010011111010000000000000000000000000000000000000000000000";
    type_cast_2221_wire_constant <= "0100000010100011100010000000000000000000000000000000000000000000";
    type_cast_2234_wire_constant <= "10111001010100011011011100010111";
    type_cast_2240_wire_constant <= "00111111101100110011001100110011";
    type_cast_2246_wire_constant <= "01000011100101100000000000000000";
    type_cast_2254_wire_constant <= "0100000010100111011100000000000000000000000000000000000000000000";
    type_cast_2267_wire_constant <= "10111001101111001011111001100010";
    type_cast_2273_wire_constant <= "00111111111001100110011001100110";
    type_cast_2279_wire_constant <= "01000011100101100000000000000000";
    type_cast_2287_wire_constant <= "10111001110111000011001101110010";
    type_cast_2293_wire_constant <= "00111111111111010111000010100100";
    type_cast_2299_wire_constant <= "01000011100101100000000000000000";
    type_cast_2314_wire_constant <= "01000011100101100000000000000000";
    type_cast_2319_wire_constant <= "01000010001000011110101110000101";
    type_cast_2325_wire_constant <= "01000010110011111101011011110000";
    type_cast_2340_wire_constant <= "00000000000000000000000000000000";
    type_cast_2353_wire_constant <= "00000000000000000000000000000111";
    type_cast_2359_wire_constant <= "00111111111111111111111110000000";
    type_cast_2365_wire_constant <= "01000000000000000000000000000000";
    type_cast_2382_wire_constant <= "00000000000000000000000000000000";
    type_cast_2387_wire_constant <= "00000000000000000000000000000001";
    type_cast_2393_wire_constant <= "00000000000000011001111111100001";
    type_cast_2411_wire_constant <= "00000000000000011001111111100001";
    type_cast_2418_wire_constant <= "00000000000000000000000000000001";
    type_cast_2423_wire_constant <= "00000000000000000000000000000001";
    type_cast_2429_wire_constant <= "00000000000000000000000000000001";
    type_cast_2459_wire_constant <= "00000000000000011001111111100001";
    type_cast_2466_wire_constant <= "00000000000000000000000000000001";
    type_cast_2483_wire_constant <= "00000000000000011001111111100001";
    type_cast_2501_wire_constant <= "00000000000000000000000000010111";
    type_cast_2507_wire_constant <= "10000000000000000000000000000000";
    type_cast_2513_wire_constant <= "00000000000000000000000011111111";
    type_cast_2519_wire_constant <= "11111111111111111111111101111011";
    type_cast_2525_wire_constant <= "00000000100000000000000000000000";
    type_cast_2531_wire_constant <= "00000000000000000000000000000000";
    type_cast_2539_wire_constant <= "00000000000000000000000000000000";
    type_cast_2562_wire_constant <= "00000000000000000000000000000000";
    type_cast_2573_wire_constant <= "00000000000000000000000000000001";
    type_cast_2579_wire_constant <= "00000000100000000000000000000000";
    type_cast_2585_wire_constant <= "00000000000000000000000000000000";
    type_cast_2593_wire_constant <= "00000000000000000000000000000000";
    type_cast_2604_wire_constant <= "00000000000000000000000000000001";
    type_cast_2626_wire_constant <= "11111111111111111111111101111010";
    type_cast_2652_wire_constant <= "00000000011111111111111111111111";
    type_cast_2658_wire_constant <= "00000000000000000000000000010111";
    type_cast_2664_wire_constant <= "01000100000000000000000000000000";
    type_cast_2689_wire_constant <= "00000000000000000000000000000000";
    type_cast_2694_wire_constant <= "00111111010011110100000111110010";
    type_cast_2700_wire_constant <= "00111101110101001101001111100111";
    type_cast_2714_wire_constant <= "00000000000000000000000000000000";
    type_cast_2727_wire_constant <= "00000000000000000000000000010111";
    type_cast_2733_wire_constant <= "00000000000000000000000011111111";
    type_cast_2739_wire_constant <= "00000000000000000000000000010111";
    type_cast_2745_wire_constant <= "00000000000000000000000011111111";
    type_cast_2751_wire_constant <= "00000000000000000000000000000111";
    type_cast_2757_wire_constant <= "00111111111111111111111110000000";
    type_cast_2763_wire_constant <= "01000000000000000000000000000000";
    type_cast_2769_wire_constant <= "00000000000000000000000000000111";
    type_cast_2775_wire_constant <= "00000000000000001111111111111111";
    type_cast_2781_wire_constant <= "00000000000000010000000000000000";
    type_cast_2792_wire_constant <= "10000000000000000000000000000000";
    type_cast_2825_wire_constant <= "00000000000000000000000000000000";
    type_cast_2830_wire_constant <= "00000000000000000000000000000001";
    type_cast_2859_wire_constant <= "00000000000000000000000000000001";
    type_cast_2864_wire_constant <= "00000000000000000000000000000001";
    type_cast_2870_wire_constant <= "00000000000000000000000000000001";
    type_cast_2906_wire_constant <= "00000000000000000000000000000001";
    type_cast_2943_wire_constant <= "11111111111111111111111111111111";
    type_cast_2959_wire_constant <= "00000000100000000000000000000000";
    type_cast_2965_wire_constant <= "00000000000000000000000000000000";
    type_cast_2973_wire_constant <= "00000000000000000000000000000000";
    type_cast_2996_wire_constant <= "00000000000000000000000000000000";
    type_cast_3007_wire_constant <= "00000000000000000000000000000001";
    type_cast_3013_wire_constant <= "00000000100000000000000000000000";
    type_cast_3019_wire_constant <= "00000000000000000000000000000000";
    type_cast_3027_wire_constant <= "00000000000000000000000000000000";
    type_cast_3038_wire_constant <= "00000000000000000000000000000001";
    type_cast_3060_wire_constant <= "11111111111111111111111111111111";
    type_cast_3091_wire_constant <= "00000000011111111111111111111111";
    type_cast_3097_wire_constant <= "00000000000000000000000000010111";
    type_cast_3103_wire_constant <= "01000100000000000000000000000000";
    type_cast_3128_wire_constant <= "00000000000000000000000000000000";
    type_cast_3133_wire_constant <= "00111111100000000000000000000000";
    type_cast_3139_wire_constant <= "01000001000110110111000101110110";
    type_cast_3153_wire_constant <= "01000001000110110111000101110110";
    type_cast_3160_wire_constant <= "00000000000000000000000000000000";
    type_cast_3173_wire_constant <= "00000000000000000000000000010111";
    type_cast_3179_wire_constant <= "00000000000000000000000011111111";
    type_cast_3185_wire_constant <= "00000000000000000000000000010111";
    type_cast_3191_wire_constant <= "00000000000000000000000011111111";
    type_cast_3197_wire_constant <= "00000000000000000000000000000111";
    type_cast_3203_wire_constant <= "00111111111111111111111110000000";
    type_cast_3209_wire_constant <= "01000000000000000000000000000000";
    type_cast_3215_wire_constant <= "00000000000000000000000000000111";
    type_cast_3221_wire_constant <= "00000000000000001111111111111111";
    type_cast_3227_wire_constant <= "00000000000000010000000000000000";
    type_cast_3238_wire_constant <= "10000000000000000000000000000000";
    type_cast_3271_wire_constant <= "00000000000000000000000000000000";
    type_cast_3276_wire_constant <= "00000000000000000000000000000001";
    type_cast_3305_wire_constant <= "00000000000000000000000000000001";
    type_cast_3310_wire_constant <= "00000000000000000000000000000001";
    type_cast_3316_wire_constant <= "00000000000000000000000000000001";
    type_cast_3352_wire_constant <= "00000000000000000000000000000001";
    type_cast_3389_wire_constant <= "11111111111111111111111111111111";
    type_cast_3405_wire_constant <= "00000000100000000000000000000000";
    type_cast_3411_wire_constant <= "00000000000000000000000000000000";
    type_cast_3419_wire_constant <= "00000000000000000000000000000000";
    type_cast_3442_wire_constant <= "00000000000000000000000000000000";
    type_cast_3453_wire_constant <= "00000000000000000000000000000001";
    type_cast_3459_wire_constant <= "00000000100000000000000000000000";
    type_cast_3465_wire_constant <= "00000000000000000000000000000000";
    type_cast_3473_wire_constant <= "00000000000000000000000000000000";
    type_cast_3484_wire_constant <= "00000000000000000000000000000001";
    type_cast_3506_wire_constant <= "11111111111111111111111111111111";
    type_cast_3537_wire_constant <= "00000000011111111111111111111111";
    type_cast_3543_wire_constant <= "00000000000000000000000000010111";
    type_cast_3549_wire_constant <= "01000100000000000000000000000000";
    type_cast_3574_wire_constant <= "00000000000000000000000000000000";
    type_cast_3584_wire_constant <= "00110011010101101011111110010101";
    type_cast_3595_wire_constant <= "01000101100111000100000000000000";
    type_cast_3601_wire_constant <= "11000010110010000000000000000000";
    type_cast_3614_wire_constant <= "01000010110010000000000000000000";
    type_cast_3632_wire_constant <= "11000010110010000000000000000000";
    type_cast_3635_wire_constant <= "01000010110010000000000000000000";
    type_cast_3640_wire_constant <= "01000101011110100000000000000000";
    type_cast_3651_wire_constant <= "11000011010010000000000000000000";
    type_cast_3664_wire_constant <= "01000011010010000000000000000000";
    type_cast_3677_wire_constant <= "00000000000000000000000000000000";
    type_cast_3693_wire_constant <= "11000011010010000000000000000000";
    type_cast_3696_wire_constant <= "01000011010010000000000000000000";
    type_cast_3705_wire_constant <= "00000000000000000000000000000111";
    type_cast_3711_wire_constant <= "00111111111111111111111110000000";
    type_cast_3717_wire_constant <= "01000000000000000000000000000000";
    type_cast_3734_wire_constant <= "00000000000000000000000000000000";
    type_cast_3739_wire_constant <= "00000000000000000000000000000001";
    type_cast_3745_wire_constant <= "00000000000000010100001111010111";
    type_cast_3763_wire_constant <= "00000000000000010100001111010111";
    type_cast_3770_wire_constant <= "00000000000000000000000000000001";
    type_cast_3775_wire_constant <= "00000000000000000000000000000001";
    type_cast_3781_wire_constant <= "00000000000000000000000000000001";
    type_cast_3811_wire_constant <= "00000000000000010100001111010111";
    type_cast_3818_wire_constant <= "00000000000000000000000000000001";
    type_cast_3835_wire_constant <= "00000000000000010100001111010111";
    type_cast_3853_wire_constant <= "00000000000000000000000000010111";
    type_cast_3859_wire_constant <= "10000000000000000000000000000000";
    type_cast_3865_wire_constant <= "00000000000000000000000011111111";
    type_cast_3871_wire_constant <= "11111111111111111111111101111011";
    type_cast_3877_wire_constant <= "00000000100000000000000000000000";
    type_cast_3883_wire_constant <= "00000000000000000000000000000000";
    type_cast_3891_wire_constant <= "00000000000000000000000000000000";
    type_cast_3914_wire_constant <= "00000000000000000000000000000000";
    type_cast_3925_wire_constant <= "00000000000000000000000000000001";
    type_cast_3931_wire_constant <= "00000000100000000000000000000000";
    type_cast_3937_wire_constant <= "00000000000000000000000000000000";
    type_cast_3945_wire_constant <= "00000000000000000000000000000000";
    type_cast_3956_wire_constant <= "00000000000000000000000000000001";
    type_cast_3978_wire_constant <= "11111111111111111111111101111010";
    type_cast_4004_wire_constant <= "00000000011111111111111111111111";
    type_cast_4010_wire_constant <= "00000000000000000000000000010111";
    type_cast_4016_wire_constant <= "01000100000000000000000000000000";
    type_cast_4041_wire_constant <= "00000000000000000000000000000000";
    phi_stmt_2045: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2049_wire_constant & type_cast_2051_wire;
      req <= phi_stmt_2045_req_0 & phi_stmt_2045_req_1;
      phi: PhiBase -- 
        generic map( -- 
          num_reqs => 2,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2045_ack_0,
          idata => idata,
          odata => flux_rotor_prevx_x0_2045,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2045
    phi_stmt_2052: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2056_wire_constant & type_cast_2058_wire;
      req <= phi_stmt_2052_req_0 & phi_stmt_2052_req_1;
      phi: PhiBase -- 
        generic map( -- 
          num_reqs => 2,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2052_ack_0,
          idata => idata,
          odata => int_flux_errx_x0_2052,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2052
    phi_stmt_2059: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2063_wire_constant & type_cast_2065_wire;
      req <= phi_stmt_2059_req_0 & phi_stmt_2059_req_1;
      phi: PhiBase -- 
        generic map( -- 
          num_reqs => 2,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2059_ack_0,
          idata => idata,
          odata => int_speed_errx_x0_2059,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2059
    phi_stmt_2134: Block -- phi operator 
      signal idata: std_logic_vector(95 downto 0);
      signal req: BooleanArray(2 downto 0);
      --
    begin -- 
      idata <= type_cast_2137_wire & type_cast_2140_wire_constant & type_cast_2143_wire_constant;
      req <= phi_stmt_2134_req_0 & phi_stmt_2134_req_1 & phi_stmt_2134_req_2;
      phi: PhiBase -- 
        generic map( -- 
          num_reqs => 3,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2134_ack_0,
          idata => idata,
          odata => int_speed_errx_x1_2134,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2134
    phi_stmt_2190: Block -- phi operator 
      signal idata: std_logic_vector(95 downto 0);
      signal req: BooleanArray(2 downto 0);
      --
    begin -- 
      idata <= type_cast_2193_wire & type_cast_2196_wire_constant & type_cast_2199_wire_constant;
      req <= phi_stmt_2190_req_0 & phi_stmt_2190_req_1 & phi_stmt_2190_req_2;
      phi: PhiBase -- 
        generic map( -- 
          num_reqs => 3,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2190_ack_0,
          idata => idata,
          odata => torque_refx_x0_2190,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2190
    phi_stmt_2304: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(3 downto 0);
      --
    begin -- 
      idata <= type_cast_2307_wire & type_cast_2309_wire & type_cast_2311_wire & type_cast_2314_wire_constant;
      req <= phi_stmt_2304_req_0 & phi_stmt_2304_req_1 & phi_stmt_2304_req_2 & phi_stmt_2304_req_3;
      phi: PhiBase -- 
        generic map( -- 
          num_reqs => 4,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2304_ack_0,
          idata => idata,
          odata => flux_refx_x0_2304,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2304
    phi_stmt_2370: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2373_wire & type_cast_2375_wire;
      req <= phi_stmt_2370_req_0 & phi_stmt_2370_req_1;
      phi: PhiBase -- 
        generic map( -- 
          num_reqs => 2,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2370_ack_0,
          idata => idata,
          odata => xx_x016x_xix_xix_xi31_2370,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2370
    phi_stmt_2376: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2379_wire & type_cast_2382_wire_constant;
      req <= phi_stmt_2376_req_0 & phi_stmt_2376_req_1;
      phi: PhiBase -- 
        generic map( -- 
          num_reqs => 2,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2376_ack_0,
          idata => idata,
          odata => quotientx_x05x_xix_xix_xi32_2376,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2376
    phi_stmt_2405: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2408_wire & type_cast_2411_wire_constant;
      req <= phi_stmt_2405_req_0 & phi_stmt_2405_req_1;
      phi: PhiBase -- 
        generic map( -- 
          num_reqs => 2,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2405_ack_0,
          idata => idata,
          odata => shifted_divisorx_x03x_xix_xix_xi34_2405,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2405
    phi_stmt_2412: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2415_wire & type_cast_2418_wire_constant;
      req <= phi_stmt_2412_req_0 & phi_stmt_2412_req_1;
      phi: PhiBase -- 
        generic map( -- 
          num_reqs => 2,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2412_ack_0,
          idata => idata,
          odata => curr_quotientx_x02x_xix_xix_xi35_2412,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2412
    phi_stmt_2444: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(0 downto 0);
      --
    begin -- 
      idata <= type_cast_2447_wire;
      req(0) <= phi_stmt_2444_req_0;
      phi: PhiBase -- 
        generic map( -- 
          num_reqs => 1,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2444_ack_0,
          idata => idata,
          odata => xx_xlcssa18_2444,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2444
    phi_stmt_2448: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(0 downto 0);
      --
    begin -- 
      idata <= type_cast_2451_wire;
      req(0) <= phi_stmt_2448_req_0;
      phi: PhiBase -- 
        generic map( -- 
          num_reqs => 1,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2448_ack_0,
          idata => idata,
          odata => xx_xlcssa17_2448,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2448
    phi_stmt_2455: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2459_wire_constant & type_cast_2461_wire;
      req <= phi_stmt_2455_req_0 & phi_stmt_2455_req_1;
      phi: PhiBase -- 
        generic map( -- 
          num_reqs => 2,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2455_ack_0,
          idata => idata,
          odata => shifted_divisorx_x0x_xlcssax_xix_xix_xi37_2455,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2455
    phi_stmt_2462: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2466_wire_constant & type_cast_2468_wire;
      req <= phi_stmt_2462_req_0 & phi_stmt_2462_req_1;
      phi: PhiBase -- 
        generic map( -- 
          num_reqs => 2,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2462_ack_0,
          idata => idata,
          odata => curr_quotientx_x0x_xlcssax_xix_xix_xi38_2462,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2462
    phi_stmt_2493: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(0 downto 0);
      --
    begin -- 
      idata <= type_cast_2496_wire;
      req(0) <= phi_stmt_2493_req_0;
      phi: PhiBase -- 
        generic map( -- 
          num_reqs => 1,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2493_ack_0,
          idata => idata,
          odata => xx_xlcssa19_2493,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2493
    phi_stmt_2556: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2559_wire & type_cast_2562_wire_constant;
      req <= phi_stmt_2556_req_0 & phi_stmt_2556_req_1;
      phi: PhiBase -- 
        generic map( -- 
          num_reqs => 2,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2556_ack_0,
          idata => idata,
          odata => iNsTr_205_2556,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2556
    phi_stmt_2563: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2566_wire & type_cast_2568_wire;
      req <= phi_stmt_2563_req_0 & phi_stmt_2563_req_1;
      phi: PhiBase -- 
        generic map( -- 
          num_reqs => 2,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2563_ack_0,
          idata => idata,
          odata => tempx_x012x_xix_xi42_2563,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2563
    phi_stmt_2614: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(0 downto 0);
      --
    begin -- 
      idata <= type_cast_2617_wire;
      req(0) <= phi_stmt_2614_req_0;
      phi: PhiBase -- 
        generic map( -- 
          num_reqs => 1,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2614_ack_0,
          idata => idata,
          odata => xx_xlcssa16_2614,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2614
    phi_stmt_2618: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(0 downto 0);
      --
    begin -- 
      idata <= type_cast_2621_wire;
      req(0) <= phi_stmt_2618_req_0;
      phi: PhiBase -- 
        generic map( -- 
          num_reqs => 1,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2618_ack_0,
          idata => idata,
          odata => xx_xlcssa15_2618,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2618
    phi_stmt_2636: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2639_wire & type_cast_2641_wire;
      req <= phi_stmt_2636_req_0 & phi_stmt_2636_req_1;
      phi: PhiBase -- 
        generic map( -- 
          num_reqs => 2,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2636_ack_0,
          idata => idata,
          odata => expx_x0x_xlcssax_xix_xi49_2636,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2636
    phi_stmt_2642: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2645_wire & type_cast_2647_wire;
      req <= phi_stmt_2642_req_0 & phi_stmt_2642_req_1;
      phi: PhiBase -- 
        generic map( -- 
          num_reqs => 2,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2642_ack_0,
          idata => idata,
          odata => tempx_x0x_xlcssax_xix_xi50_2642,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2642
    phi_stmt_2683: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2686_wire & type_cast_2689_wire_constant;
      req <= phi_stmt_2683_req_0 & phi_stmt_2683_req_1;
      phi: PhiBase -- 
        generic map( -- 
          num_reqs => 2,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2683_ack_0,
          idata => idata,
          odata => iNsTr_42_2683,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2683
    phi_stmt_2813: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2816_wire & type_cast_2818_wire;
      req <= phi_stmt_2813_req_0 & phi_stmt_2813_req_1;
      phi: PhiBase -- 
        generic map( -- 
          num_reqs => 2,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2813_ack_0,
          idata => idata,
          odata => xx_x016x_xix_xix_xi3_2813,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2813
    phi_stmt_2819: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2822_wire & type_cast_2825_wire_constant;
      req <= phi_stmt_2819_req_0 & phi_stmt_2819_req_1;
      phi: PhiBase -- 
        generic map( -- 
          num_reqs => 2,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2819_ack_0,
          idata => idata,
          odata => quotientx_x05x_xix_xix_xi4_2819,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2819
    phi_stmt_2847: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2850_wire & type_cast_2852_wire;
      req <= phi_stmt_2847_req_0 & phi_stmt_2847_req_1;
      phi: PhiBase -- 
        generic map( -- 
          num_reqs => 2,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2847_ack_0,
          idata => idata,
          odata => shifted_divisorx_x03x_xix_xix_xi6_2847,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2847
    phi_stmt_2853: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2856_wire & type_cast_2859_wire_constant;
      req <= phi_stmt_2853_req_0 & phi_stmt_2853_req_1;
      phi: PhiBase -- 
        generic map( -- 
          num_reqs => 2,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2853_ack_0,
          idata => idata,
          odata => curr_quotientx_x02x_xix_xix_xi7_2853,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2853
    phi_stmt_2885: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(0 downto 0);
      --
    begin -- 
      idata <= type_cast_2888_wire;
      req(0) <= phi_stmt_2885_req_0;
      phi: PhiBase -- 
        generic map( -- 
          num_reqs => 1,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2885_ack_0,
          idata => idata,
          odata => xx_xlcssa13_2885,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2885
    phi_stmt_2889: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(0 downto 0);
      --
    begin -- 
      idata <= type_cast_2892_wire;
      req(0) <= phi_stmt_2889_req_0;
      phi: PhiBase -- 
        generic map( -- 
          num_reqs => 1,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2889_ack_0,
          idata => idata,
          odata => xx_xlcssa12_2889,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2889
    phi_stmt_2896: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2899_wire & type_cast_2901_wire;
      req <= phi_stmt_2896_req_0 & phi_stmt_2896_req_1;
      phi: PhiBase -- 
        generic map( -- 
          num_reqs => 2,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2896_ack_0,
          idata => idata,
          odata => shifted_divisorx_x0x_xlcssax_xix_xix_xi9_2896,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2896
    phi_stmt_2902: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2906_wire_constant & type_cast_2908_wire;
      req <= phi_stmt_2902_req_0 & phi_stmt_2902_req_1;
      phi: PhiBase -- 
        generic map( -- 
          num_reqs => 2,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2902_ack_0,
          idata => idata,
          odata => curr_quotientx_x0x_xlcssax_xix_xix_xi10_2902,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2902
    phi_stmt_2932: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(0 downto 0);
      --
    begin -- 
      idata <= type_cast_2935_wire;
      req(0) <= phi_stmt_2932_req_0;
      phi: PhiBase -- 
        generic map( -- 
          num_reqs => 1,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2932_ack_0,
          idata => idata,
          odata => xx_xlcssa14_2932,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2932
    phi_stmt_2939: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2943_wire_constant & type_cast_2945_wire;
      req <= phi_stmt_2939_req_0 & phi_stmt_2939_req_1;
      phi: PhiBase -- 
        generic map( -- 
          num_reqs => 2,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2939_ack_0,
          idata => idata,
          odata => xx_x0x_xix_xix_xi12_2939,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2939
    phi_stmt_2949: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2952_wire & type_cast_2954_wire;
      req <= phi_stmt_2949_req_0 & phi_stmt_2949_req_1;
      phi: PhiBase -- 
        generic map( -- 
          num_reqs => 2,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2949_ack_0,
          idata => idata,
          odata => tempx_x0x_xphx_xix_xi14_2949,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2949
    phi_stmt_2990: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2993_wire & type_cast_2996_wire_constant;
      req <= phi_stmt_2990_req_0 & phi_stmt_2990_req_1;
      phi: PhiBase -- 
        generic map( -- 
          num_reqs => 2,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2990_ack_0,
          idata => idata,
          odata => iNsTr_169_2990,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2990
    phi_stmt_2997: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_3000_wire & type_cast_3002_wire;
      req <= phi_stmt_2997_req_0 & phi_stmt_2997_req_1;
      phi: PhiBase -- 
        generic map( -- 
          num_reqs => 2,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2997_ack_0,
          idata => idata,
          odata => tempx_x012x_xix_xi17_2997,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2997
    phi_stmt_3048: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(0 downto 0);
      --
    begin -- 
      idata <= type_cast_3051_wire;
      req(0) <= phi_stmt_3048_req_0;
      phi: PhiBase -- 
        generic map( -- 
          num_reqs => 1,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_3048_ack_0,
          idata => idata,
          odata => xx_xlcssa11_3048,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_3048
    phi_stmt_3052: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(0 downto 0);
      --
    begin -- 
      idata <= type_cast_3055_wire;
      req(0) <= phi_stmt_3052_req_0;
      phi: PhiBase -- 
        generic map( -- 
          num_reqs => 1,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_3052_ack_0,
          idata => idata,
          odata => xx_xlcssa10_3052,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_3052
    phi_stmt_3075: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_3078_wire & type_cast_3080_wire;
      req <= phi_stmt_3075_req_0 & phi_stmt_3075_req_1;
      phi: PhiBase -- 
        generic map( -- 
          num_reqs => 2,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_3075_ack_0,
          idata => idata,
          odata => expx_x0x_xlcssax_xix_xi25_3075,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_3075
    phi_stmt_3081: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_3084_wire & type_cast_3086_wire;
      req <= phi_stmt_3081_req_0 & phi_stmt_3081_req_1;
      phi: PhiBase -- 
        generic map( -- 
          num_reqs => 2,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_3081_ack_0,
          idata => idata,
          odata => tempx_x0x_xlcssax_xix_xi26_3081,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_3081
    phi_stmt_3122: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_3125_wire & type_cast_3128_wire_constant;
      req <= phi_stmt_3122_req_0 & phi_stmt_3122_req_1;
      phi: PhiBase -- 
        generic map( -- 
          num_reqs => 2,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_3122_ack_0,
          idata => idata,
          odata => iNsTr_59_3122,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_3122
    phi_stmt_3259: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_3262_wire & type_cast_3264_wire;
      req <= phi_stmt_3259_req_0 & phi_stmt_3259_req_1;
      phi: PhiBase -- 
        generic map( -- 
          num_reqs => 2,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_3259_ack_0,
          idata => idata,
          odata => xx_x016x_xix_xix_xi_3259,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_3259
    phi_stmt_3265: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_3268_wire & type_cast_3271_wire_constant;
      req <= phi_stmt_3265_req_0 & phi_stmt_3265_req_1;
      phi: PhiBase -- 
        generic map( -- 
          num_reqs => 2,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_3265_ack_0,
          idata => idata,
          odata => quotientx_x05x_xix_xix_xi_3265,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_3265
    phi_stmt_3293: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_3296_wire & type_cast_3298_wire;
      req <= phi_stmt_3293_req_0 & phi_stmt_3293_req_1;
      phi: PhiBase -- 
        generic map( -- 
          num_reqs => 2,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_3293_ack_0,
          idata => idata,
          odata => shifted_divisorx_x03x_xix_xix_xi_3293,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_3293
    phi_stmt_3299: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_3302_wire & type_cast_3305_wire_constant;
      req <= phi_stmt_3299_req_0 & phi_stmt_3299_req_1;
      phi: PhiBase -- 
        generic map( -- 
          num_reqs => 2,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_3299_ack_0,
          idata => idata,
          odata => curr_quotientx_x02x_xix_xix_xi_3299,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_3299
    phi_stmt_3331: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(0 downto 0);
      --
    begin -- 
      idata <= type_cast_3334_wire;
      req(0) <= phi_stmt_3331_req_0;
      phi: PhiBase -- 
        generic map( -- 
          num_reqs => 1,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_3331_ack_0,
          idata => idata,
          odata => xx_xlcssa8_3331,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_3331
    phi_stmt_3335: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(0 downto 0);
      --
    begin -- 
      idata <= type_cast_3338_wire;
      req(0) <= phi_stmt_3335_req_0;
      phi: PhiBase -- 
        generic map( -- 
          num_reqs => 1,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_3335_ack_0,
          idata => idata,
          odata => xx_xlcssa7_3335,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_3335
    phi_stmt_3342: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_3345_wire & type_cast_3347_wire;
      req <= phi_stmt_3342_req_0 & phi_stmt_3342_req_1;
      phi: PhiBase -- 
        generic map( -- 
          num_reqs => 2,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_3342_ack_0,
          idata => idata,
          odata => shifted_divisorx_x0x_xlcssax_xix_xix_xi_3342,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_3342
    phi_stmt_3348: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_3352_wire_constant & type_cast_3354_wire;
      req <= phi_stmt_3348_req_0 & phi_stmt_3348_req_1;
      phi: PhiBase -- 
        generic map( -- 
          num_reqs => 2,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_3348_ack_0,
          idata => idata,
          odata => curr_quotientx_x0x_xlcssax_xix_xix_xi_3348,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_3348
    phi_stmt_3378: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(0 downto 0);
      --
    begin -- 
      idata <= type_cast_3381_wire;
      req(0) <= phi_stmt_3378_req_0;
      phi: PhiBase -- 
        generic map( -- 
          num_reqs => 1,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_3378_ack_0,
          idata => idata,
          odata => xx_xlcssa9_3378,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_3378
    phi_stmt_3385: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_3389_wire_constant & type_cast_3391_wire;
      req <= phi_stmt_3385_req_0 & phi_stmt_3385_req_1;
      phi: PhiBase -- 
        generic map( -- 
          num_reqs => 2,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_3385_ack_0,
          idata => idata,
          odata => xx_x0x_xix_xix_xi_3385,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_3385
    phi_stmt_3395: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_3398_wire & type_cast_3400_wire;
      req <= phi_stmt_3395_req_0 & phi_stmt_3395_req_1;
      phi: PhiBase -- 
        generic map( -- 
          num_reqs => 2,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_3395_ack_0,
          idata => idata,
          odata => tempx_x0x_xphx_xix_xi_3395,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_3395
    phi_stmt_3436: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_3439_wire & type_cast_3442_wire_constant;
      req <= phi_stmt_3436_req_0 & phi_stmt_3436_req_1;
      phi: PhiBase -- 
        generic map( -- 
          num_reqs => 2,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_3436_ack_0,
          idata => idata,
          odata => iNsTr_193_3436,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_3436
    phi_stmt_3443: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_3446_wire & type_cast_3448_wire;
      req <= phi_stmt_3443_req_0 & phi_stmt_3443_req_1;
      phi: PhiBase -- 
        generic map( -- 
          num_reqs => 2,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_3443_ack_0,
          idata => idata,
          odata => tempx_x012x_xix_xi_3443,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_3443
    phi_stmt_3494: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(0 downto 0);
      --
    begin -- 
      idata <= type_cast_3497_wire;
      req(0) <= phi_stmt_3494_req_0;
      phi: PhiBase -- 
        generic map( -- 
          num_reqs => 1,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_3494_ack_0,
          idata => idata,
          odata => xx_xlcssa6_3494,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_3494
    phi_stmt_3498: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(0 downto 0);
      --
    begin -- 
      idata <= type_cast_3501_wire;
      req(0) <= phi_stmt_3498_req_0;
      phi: PhiBase -- 
        generic map( -- 
          num_reqs => 1,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_3498_ack_0,
          idata => idata,
          odata => xx_xlcssa5_3498,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_3498
    phi_stmt_3521: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_3524_wire & type_cast_3526_wire;
      req <= phi_stmt_3521_req_0 & phi_stmt_3521_req_1;
      phi: PhiBase -- 
        generic map( -- 
          num_reqs => 2,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_3521_ack_0,
          idata => idata,
          odata => expx_x0x_xlcssax_xix_xi_3521,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_3521
    phi_stmt_3527: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_3530_wire & type_cast_3532_wire;
      req <= phi_stmt_3527_req_0 & phi_stmt_3527_req_1;
      phi: PhiBase -- 
        generic map( -- 
          num_reqs => 2,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_3527_ack_0,
          idata => idata,
          odata => tempx_x0x_xlcssax_xix_xi_3527,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_3527
    phi_stmt_3568: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_3571_wire & type_cast_3574_wire_constant;
      req <= phi_stmt_3568_req_0 & phi_stmt_3568_req_1;
      phi: PhiBase -- 
        generic map( -- 
          num_reqs => 2,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_3568_ack_0,
          idata => idata,
          odata => iNsTr_81_3568,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_3568
    phi_stmt_3626: Block -- phi operator 
      signal idata: std_logic_vector(95 downto 0);
      signal req: BooleanArray(2 downto 0);
      --
    begin -- 
      idata <= type_cast_3629_wire & type_cast_3632_wire_constant & type_cast_3635_wire_constant;
      req <= phi_stmt_3626_req_0 & phi_stmt_3626_req_1 & phi_stmt_3626_req_2;
      phi: PhiBase -- 
        generic map( -- 
          num_reqs => 3,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_3626_ack_0,
          idata => idata,
          odata => int_flux_errx_x1_3626,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_3626
    phi_stmt_3687: Block -- phi operator 
      signal idata: std_logic_vector(95 downto 0);
      signal req: BooleanArray(2 downto 0);
      --
    begin -- 
      idata <= type_cast_3690_wire & type_cast_3693_wire_constant & type_cast_3696_wire_constant;
      req <= phi_stmt_3687_req_0 & phi_stmt_3687_req_1 & phi_stmt_3687_req_2;
      phi: PhiBase -- 
        generic map( -- 
          num_reqs => 3,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_3687_ack_0,
          idata => idata,
          odata => tmp10x_xi55x_xin_3687,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_3687
    phi_stmt_3722: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_3725_wire & type_cast_3727_wire;
      req <= phi_stmt_3722_req_0 & phi_stmt_3722_req_1;
      phi: PhiBase -- 
        generic map( -- 
          num_reqs => 2,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_3722_ack_0,
          idata => idata,
          odata => xx_x016x_xix_xi_3722,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_3722
    phi_stmt_3728: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_3731_wire & type_cast_3734_wire_constant;
      req <= phi_stmt_3728_req_0 & phi_stmt_3728_req_1;
      phi: PhiBase -- 
        generic map( -- 
          num_reqs => 2,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_3728_ack_0,
          idata => idata,
          odata => quotientx_x05x_xix_xi_3728,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_3728
    phi_stmt_3757: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_3760_wire & type_cast_3763_wire_constant;
      req <= phi_stmt_3757_req_0 & phi_stmt_3757_req_1;
      phi: PhiBase -- 
        generic map( -- 
          num_reqs => 2,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_3757_ack_0,
          idata => idata,
          odata => shifted_divisorx_x03x_xix_xi_3757,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_3757
    phi_stmt_3764: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_3767_wire & type_cast_3770_wire_constant;
      req <= phi_stmt_3764_req_0 & phi_stmt_3764_req_1;
      phi: PhiBase -- 
        generic map( -- 
          num_reqs => 2,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_3764_ack_0,
          idata => idata,
          odata => curr_quotientx_x02x_xix_xi_3764,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_3764
    phi_stmt_3796: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(0 downto 0);
      --
    begin -- 
      idata <= type_cast_3799_wire;
      req(0) <= phi_stmt_3796_req_0;
      phi: PhiBase -- 
        generic map( -- 
          num_reqs => 1,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_3796_ack_0,
          idata => idata,
          odata => xx_xlcssa3_3796,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_3796
    phi_stmt_3800: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(0 downto 0);
      --
    begin -- 
      idata <= type_cast_3803_wire;
      req(0) <= phi_stmt_3800_req_0;
      phi: PhiBase -- 
        generic map( -- 
          num_reqs => 1,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_3800_ack_0,
          idata => idata,
          odata => xx_xlcssa2_3800,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_3800
    phi_stmt_3807: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_3811_wire_constant & type_cast_3813_wire;
      req <= phi_stmt_3807_req_0 & phi_stmt_3807_req_1;
      phi: PhiBase -- 
        generic map( -- 
          num_reqs => 2,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_3807_ack_0,
          idata => idata,
          odata => shifted_divisorx_x0x_xlcssax_xix_xi_3807,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_3807
    phi_stmt_3814: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_3818_wire_constant & type_cast_3820_wire;
      req <= phi_stmt_3814_req_0 & phi_stmt_3814_req_1;
      phi: PhiBase -- 
        generic map( -- 
          num_reqs => 2,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_3814_ack_0,
          idata => idata,
          odata => curr_quotientx_x0x_xlcssax_xix_xi_3814,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_3814
    phi_stmt_3845: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(0 downto 0);
      --
    begin -- 
      idata <= type_cast_3848_wire;
      req(0) <= phi_stmt_3845_req_0;
      phi: PhiBase -- 
        generic map( -- 
          num_reqs => 1,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_3845_ack_0,
          idata => idata,
          odata => xx_xlcssa4_3845,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_3845
    phi_stmt_3908: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_3911_wire & type_cast_3914_wire_constant;
      req <= phi_stmt_3908_req_0 & phi_stmt_3908_req_1;
      phi: PhiBase -- 
        generic map( -- 
          num_reqs => 2,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_3908_ack_0,
          idata => idata,
          odata => iNsTr_255_3908,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_3908
    phi_stmt_3915: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_3918_wire & type_cast_3920_wire;
      req <= phi_stmt_3915_req_0 & phi_stmt_3915_req_1;
      phi: PhiBase -- 
        generic map( -- 
          num_reqs => 2,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_3915_ack_0,
          idata => idata,
          odata => tempx_x012x_xi_3915,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_3915
    phi_stmt_3966: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(0 downto 0);
      --
    begin -- 
      idata <= type_cast_3969_wire;
      req(0) <= phi_stmt_3966_req_0;
      phi: PhiBase -- 
        generic map( -- 
          num_reqs => 1,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_3966_ack_0,
          idata => idata,
          odata => xx_xlcssa1_3966,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_3966
    phi_stmt_3970: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(0 downto 0);
      --
    begin -- 
      idata <= type_cast_3973_wire;
      req(0) <= phi_stmt_3970_req_0;
      phi: PhiBase -- 
        generic map( -- 
          num_reqs => 1,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_3970_ack_0,
          idata => idata,
          odata => xx_xlcssa_3970,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_3970
    phi_stmt_3988: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_3991_wire & type_cast_3993_wire;
      req <= phi_stmt_3988_req_0 & phi_stmt_3988_req_1;
      phi: PhiBase -- 
        generic map( -- 
          num_reqs => 2,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_3988_ack_0,
          idata => idata,
          odata => expx_x0x_xlcssax_xi_3988,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_3988
    phi_stmt_3994: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_3997_wire & type_cast_3999_wire;
      req <= phi_stmt_3994_req_0 & phi_stmt_3994_req_1;
      phi: PhiBase -- 
        generic map( -- 
          num_reqs => 2,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_3994_ack_0,
          idata => idata,
          odata => tempx_x0x_xlcssax_xi_3994,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_3994
    phi_stmt_4035: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_4038_wire & type_cast_4041_wire_constant;
      req <= phi_stmt_4035_req_0 & phi_stmt_4035_req_1;
      phi: PhiBase -- 
        generic map( -- 
          num_reqs => 2,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_4035_ack_0,
          idata => idata,
          odata => iNsTr_216_4035,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_4035
    MUX_3155_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= MUX_3155_inst_req_0;
      MUX_3155_inst_ack_0<= sample_ack(0);
      update_req(0) <= MUX_3155_inst_req_1;
      MUX_3155_inst_ack_1<= update_ack(0);
      MUX_3155_inst: SelectSplitProtocol generic map(name => "MUX_3155_inst", data_width => 32, buffering => 1, flow_through => false) -- 
        port map( x => type_cast_3153_wire_constant, y => iNsTr_61_3149, sel => iNsTr_60_3135, z => tmp6x_xix_xi_3156, sample_req => sample_req(0), sample_ack => sample_ack(0), update_req => update_req(0), update_ack => update_ack(0), clk => clk, reset => reset); -- 
      -- 
    end block;
    type_cast_2051_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2051_inst_req_0;
      type_cast_2051_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2051_inst_req_1;
      type_cast_2051_inst_ack_1<= rack(0);
      type_cast_2051_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2051_inst",
        buffer_size => 1,
        in_data_width => 32,
        out_data_width => 32
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => iNsTr_42_2683,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2051_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2058_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2058_inst_req_0;
      type_cast_2058_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2058_inst_req_1;
      type_cast_2058_inst_ack_1<= rack(0);
      type_cast_2058_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2058_inst",
        buffer_size => 1,
        in_data_width => 32,
        out_data_width => 32
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => int_flux_errx_x1_3626,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2058_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2065_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2065_inst_req_0;
      type_cast_2065_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2065_inst_req_1;
      type_cast_2065_inst_ack_1<= rack(0);
      type_cast_2065_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2065_inst",
        buffer_size => 1,
        in_data_width => 32,
        out_data_width => 32
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => int_speed_errx_x1_2134,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2065_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2137_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2137_inst_req_0;
      type_cast_2137_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2137_inst_req_1;
      type_cast_2137_inst_ack_1<= rack(0);
      type_cast_2137_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2137_inst",
        buffer_size => 1,
        in_data_width => 32,
        out_data_width => 32
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => iNsTr_12_2100,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2137_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2193_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2193_inst_req_0;
      type_cast_2193_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2193_inst_req_1;
      type_cast_2193_inst_ack_1<= rack(0);
      type_cast_2193_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2193_inst",
        buffer_size => 1,
        in_data_width => 32,
        out_data_width => 32
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => phitmp_2187,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2193_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2307_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2307_inst_req_0;
      type_cast_2307_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2307_inst_req_1;
      type_cast_2307_inst_ack_1<= rack(0);
      type_cast_2307_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2307_inst",
        buffer_size => 1,
        in_data_width => 32,
        out_data_width => 32
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => iNsTr_40_2248,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2307_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2309_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2309_inst_req_0;
      type_cast_2309_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2309_inst_req_1;
      type_cast_2309_inst_ack_1<= rack(0);
      type_cast_2309_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2309_inst",
        buffer_size => 1,
        in_data_width => 32,
        out_data_width => 32
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => iNsTr_57_2281,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2309_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2311_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2311_inst_req_0;
      type_cast_2311_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2311_inst_req_1;
      type_cast_2311_inst_ack_1<= rack(0);
      type_cast_2311_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2311_inst",
        buffer_size => 1,
        in_data_width => 32,
        out_data_width => 32
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => iNsTr_53_2301,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2311_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2335_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2335_inst_req_0;
      type_cast_2335_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2335_inst_req_1;
      type_cast_2335_inst_ack_1<= rack(0);
      type_cast_2335_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2335_inst",
        buffer_size => 1,
        in_data_width => 32,
        out_data_width => 32
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => iNsTr_32_2332,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp10x_xix_xi30_2336,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2373_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2373_inst_req_0;
      type_cast_2373_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2373_inst_req_1;
      type_cast_2373_inst_ack_1<= rack(0);
      type_cast_2373_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2373_inst",
        buffer_size => 1,
        in_data_width => 32,
        out_data_width => 32
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => iNsTr_110_2479,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2373_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2375_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2375_inst_req_0;
      type_cast_2375_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2375_inst_req_1;
      type_cast_2375_inst_ack_1<= rack(0);
      type_cast_2375_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2375_inst",
        buffer_size => 1,
        in_data_width => 32,
        out_data_width => 32
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => iNsTr_49_2367,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2375_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2379_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2379_inst_req_0;
      type_cast_2379_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2379_inst_req_1;
      type_cast_2379_inst_ack_1<= rack(0);
      type_cast_2379_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2379_inst",
        buffer_size => 1,
        in_data_width => 32,
        out_data_width => 32
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => iNsTr_109_2474,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2379_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2408_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2408_inst_req_0;
      type_cast_2408_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2408_inst_req_1;
      type_cast_2408_inst_ack_1<= rack(0);
      type_cast_2408_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2408_inst",
        buffer_size => 1,
        in_data_width => 32,
        out_data_width => 32
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => iNsTr_135_2425,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2408_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2415_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2415_inst_req_0;
      type_cast_2415_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2415_inst_req_1;
      type_cast_2415_inst_ack_1<= rack(0);
      type_cast_2415_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2415_inst",
        buffer_size => 1,
        in_data_width => 32,
        out_data_width => 32
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => iNsTr_136_2431,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2415_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2447_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2447_inst_req_0;
      type_cast_2447_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2447_inst_req_1;
      type_cast_2447_inst_ack_1<= rack(0);
      type_cast_2447_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2447_inst",
        buffer_size => 1,
        in_data_width => 32,
        out_data_width => 32
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => iNsTr_136_2431,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2447_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2451_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2451_inst_req_0;
      type_cast_2451_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2451_inst_req_1;
      type_cast_2451_inst_ack_1<= rack(0);
      type_cast_2451_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2451_inst",
        buffer_size => 1,
        in_data_width => 32,
        out_data_width => 32
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => iNsTr_135_2425,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2451_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2461_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2461_inst_req_0;
      type_cast_2461_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2461_inst_req_1;
      type_cast_2461_inst_ack_1<= rack(0);
      type_cast_2461_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2461_inst",
        buffer_size => 1,
        in_data_width => 32,
        out_data_width => 32
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => xx_xlcssa17_2448,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2461_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2468_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2468_inst_req_0;
      type_cast_2468_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2468_inst_req_1;
      type_cast_2468_inst_ack_1<= rack(0);
      type_cast_2468_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2468_inst",
        buffer_size => 1,
        in_data_width => 32,
        out_data_width => 32
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => xx_xlcssa18_2444,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2468_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2496_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2496_inst_req_0;
      type_cast_2496_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2496_inst_req_1;
      type_cast_2496_inst_ack_1<= rack(0);
      type_cast_2496_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2496_inst",
        buffer_size => 1,
        in_data_width => 32,
        out_data_width => 32
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => iNsTr_109_2474,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2496_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2559_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2559_inst_req_0;
      type_cast_2559_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2559_inst_req_1;
      type_cast_2559_inst_ack_1<= rack(0);
      type_cast_2559_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2559_inst",
        buffer_size => 1,
        in_data_width => 32,
        out_data_width => 32
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnextx_xix_xi44_2606,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2559_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2566_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2566_inst_req_0;
      type_cast_2566_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2566_inst_req_1;
      type_cast_2566_inst_ack_1<= rack(0);
      type_cast_2566_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2566_inst",
        buffer_size => 1,
        in_data_width => 32,
        out_data_width => 32
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => iNsTr_206_2575,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2566_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2568_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2568_inst_req_0;
      type_cast_2568_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2568_inst_req_1;
      type_cast_2568_inst_ack_1<= rack(0);
      type_cast_2568_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2568_inst",
        buffer_size => 1,
        in_data_width => 32,
        out_data_width => 32
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => xx_xlcssa19_2493,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2568_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2617_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2617_inst_req_0;
      type_cast_2617_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2617_inst_req_1;
      type_cast_2617_inst_ack_1<= rack(0);
      type_cast_2617_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2617_inst",
        buffer_size => 1,
        in_data_width => 32,
        out_data_width => 32
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => iNsTr_206_2575,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2617_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2621_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2621_inst_req_0;
      type_cast_2621_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2621_inst_req_1;
      type_cast_2621_inst_ack_1<= rack(0);
      type_cast_2621_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2621_inst",
        buffer_size => 1,
        in_data_width => 32,
        out_data_width => 32
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => iNsTr_205_2556,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2621_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2639_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2639_inst_req_0;
      type_cast_2639_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2639_inst_req_1;
      type_cast_2639_inst_ack_1<= rack(0);
      type_cast_2639_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2639_inst",
        buffer_size => 1,
        in_data_width => 32,
        out_data_width => 32
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp26x_xix_xi47_2633,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2639_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2641_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2641_inst_req_0;
      type_cast_2641_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2641_inst_req_1;
      type_cast_2641_inst_ack_1<= rack(0);
      type_cast_2641_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2641_inst",
        buffer_size => 1,
        in_data_width => 32,
        out_data_width => 32
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => iNsTr_142_2521,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2641_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2645_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2645_inst_req_0;
      type_cast_2645_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2645_inst_req_1;
      type_cast_2645_inst_ack_1<= rack(0);
      type_cast_2645_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2645_inst",
        buffer_size => 1,
        in_data_width => 32,
        out_data_width => 32
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => xx_xlcssa16_2614,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2645_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2647_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2647_inst_req_0;
      type_cast_2647_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2647_inst_req_1;
      type_cast_2647_inst_ack_1<= rack(0);
      type_cast_2647_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2647_inst",
        buffer_size => 1,
        in_data_width => 32,
        out_data_width => 32
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => xx_xlcssa19_2493,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2647_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2679_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2679_inst_req_0;
      type_cast_2679_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2679_inst_req_1;
      type_cast_2679_inst_ack_1<= rack(0);
      type_cast_2679_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2679_inst",
        buffer_size => 1,
        in_data_width => 32,
        out_data_width => 32
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => iNsTr_181_2676,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp3x_xix_xi51_2680,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2686_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2686_inst_req_0;
      type_cast_2686_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2686_inst_req_1;
      type_cast_2686_inst_ack_1<= rack(0);
      type_cast_2686_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2686_inst",
        buffer_size => 1,
        in_data_width => 32,
        out_data_width => 32
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp3x_xix_xi51_2680,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2686_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2705_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2705_inst_req_0;
      type_cast_2705_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2705_inst_req_1;
      type_cast_2705_inst_ack_1<= rack(0);
      type_cast_2705_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2705_inst",
        buffer_size => 1,
        in_data_width => 32,
        out_data_width => 32
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => iNsTr_43_2696,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp10x_xix_xi1_2706,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2709_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2709_inst_req_0;
      type_cast_2709_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2709_inst_req_1;
      type_cast_2709_inst_ack_1<= rack(0);
      type_cast_2709_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2709_inst",
        buffer_size => 1,
        in_data_width => 32,
        out_data_width => 32
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => iNsTr_44_2702,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp6x_xix_xi2_2710,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2816_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2816_inst_req_0;
      type_cast_2816_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2816_inst_req_1;
      type_cast_2816_inst_ack_1<= rack(0);
      type_cast_2816_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2816_inst",
        buffer_size => 1,
        in_data_width => 32,
        out_data_width => 32
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => iNsTr_166_2919,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2816_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2818_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2818_inst_req_0;
      type_cast_2818_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2818_inst_req_1;
      type_cast_2818_inst_ack_1<= rack(0);
      type_cast_2818_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2818_inst",
        buffer_size => 1,
        in_data_width => 32,
        out_data_width => 32
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => iNsTr_70_2765,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2818_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2822_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2822_inst_req_0;
      type_cast_2822_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2822_inst_req_1;
      type_cast_2822_inst_ack_1<= rack(0);
      type_cast_2822_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2822_inst",
        buffer_size => 1,
        in_data_width => 32,
        out_data_width => 32
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => iNsTr_165_2914,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2822_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2850_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2850_inst_req_0;
      type_cast_2850_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2850_inst_req_1;
      type_cast_2850_inst_ack_1<= rack(0);
      type_cast_2850_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2850_inst",
        buffer_size => 1,
        in_data_width => 32,
        out_data_width => 32
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => iNsTr_199_2866,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2850_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2852_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2852_inst_req_0;
      type_cast_2852_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2852_inst_req_1;
      type_cast_2852_inst_ack_1<= rack(0);
      type_cast_2852_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2852_inst",
        buffer_size => 1,
        in_data_width => 32,
        out_data_width => 32
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => iNsTr_73_2783,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2852_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2856_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2856_inst_req_0;
      type_cast_2856_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2856_inst_req_1;
      type_cast_2856_inst_ack_1<= rack(0);
      type_cast_2856_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2856_inst",
        buffer_size => 1,
        in_data_width => 32,
        out_data_width => 32
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => iNsTr_200_2872,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2856_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2888_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2888_inst_req_0;
      type_cast_2888_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2888_inst_req_1;
      type_cast_2888_inst_ack_1<= rack(0);
      type_cast_2888_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2888_inst",
        buffer_size => 1,
        in_data_width => 32,
        out_data_width => 32
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => iNsTr_200_2872,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2888_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2892_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2892_inst_req_0;
      type_cast_2892_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2892_inst_req_1;
      type_cast_2892_inst_ack_1<= rack(0);
      type_cast_2892_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2892_inst",
        buffer_size => 1,
        in_data_width => 32,
        out_data_width => 32
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => iNsTr_199_2866,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2892_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2899_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2899_inst_req_0;
      type_cast_2899_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2899_inst_req_1;
      type_cast_2899_inst_ack_1<= rack(0);
      type_cast_2899_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2899_inst",
        buffer_size => 1,
        in_data_width => 32,
        out_data_width => 32
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => iNsTr_73_2783,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2899_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2901_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2901_inst_req_0;
      type_cast_2901_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2901_inst_req_1;
      type_cast_2901_inst_ack_1<= rack(0);
      type_cast_2901_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2901_inst",
        buffer_size => 1,
        in_data_width => 32,
        out_data_width => 32
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => xx_xlcssa12_2889,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2901_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2908_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2908_inst_req_0;
      type_cast_2908_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2908_inst_req_1;
      type_cast_2908_inst_ack_1<= rack(0);
      type_cast_2908_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2908_inst",
        buffer_size => 1,
        in_data_width => 32,
        out_data_width => 32
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => xx_xlcssa13_2885,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2908_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2935_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2935_inst_req_0;
      type_cast_2935_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2935_inst_req_1;
      type_cast_2935_inst_ack_1<= rack(0);
      type_cast_2935_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2935_inst",
        buffer_size => 1,
        in_data_width => 32,
        out_data_width => 32
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => iNsTr_165_2914,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2935_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2945_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2945_inst_req_0;
      type_cast_2945_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2945_inst_req_1;
      type_cast_2945_inst_ack_1<= rack(0);
      type_cast_2945_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2945_inst",
        buffer_size => 1,
        in_data_width => 32,
        out_data_width => 32
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => xx_xlcssa14_2932,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2945_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2952_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2952_inst_req_0;
      type_cast_2952_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2952_inst_req_1;
      type_cast_2952_inst_ack_1<= rack(0);
      type_cast_2952_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2952_inst",
        buffer_size => 1,
        in_data_width => 32,
        out_data_width => 32
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => xx_x0x_xix_xix_xi12_2939,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2952_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2954_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2954_inst_req_0;
      type_cast_2954_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2954_inst_req_1;
      type_cast_2954_inst_ack_1<= rack(0);
      type_cast_2954_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2954_inst",
        buffer_size => 1,
        in_data_width => 32,
        out_data_width => 32
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => iNsTr_70_2765,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2954_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2993_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2993_inst_req_0;
      type_cast_2993_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2993_inst_req_1;
      type_cast_2993_inst_ack_1<= rack(0);
      type_cast_2993_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2993_inst",
        buffer_size => 1,
        in_data_width => 32,
        out_data_width => 32
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnextx_xix_xi19_3040,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2993_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3000_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3000_inst_req_0;
      type_cast_3000_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3000_inst_req_1;
      type_cast_3000_inst_ack_1<= rack(0);
      type_cast_3000_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3000_inst",
        buffer_size => 1,
        in_data_width => 32,
        out_data_width => 32
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => iNsTr_170_3009,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_3000_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3002_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3002_inst_req_0;
      type_cast_3002_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3002_inst_req_1;
      type_cast_3002_inst_ack_1<= rack(0);
      type_cast_3002_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3002_inst",
        buffer_size => 1,
        in_data_width => 32,
        out_data_width => 32
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tempx_x0x_xphx_xix_xi14_2949,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_3002_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3051_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3051_inst_req_0;
      type_cast_3051_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3051_inst_req_1;
      type_cast_3051_inst_ack_1<= rack(0);
      type_cast_3051_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3051_inst",
        buffer_size => 1,
        in_data_width => 32,
        out_data_width => 32
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => iNsTr_170_3009,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_3051_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3055_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3055_inst_req_0;
      type_cast_3055_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3055_inst_req_1;
      type_cast_3055_inst_ack_1<= rack(0);
      type_cast_3055_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3055_inst",
        buffer_size => 1,
        in_data_width => 32,
        out_data_width => 32
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => iNsTr_169_2990,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_3055_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3078_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3078_inst_req_0;
      type_cast_3078_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3078_inst_req_1;
      type_cast_3078_inst_ack_1<= rack(0);
      type_cast_3078_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3078_inst",
        buffer_size => 1,
        in_data_width => 32,
        out_data_width => 32
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp26x_xix_xi23_3072,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_3078_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3080_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3080_inst_req_0;
      type_cast_3080_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3080_inst_req_1;
      type_cast_3080_inst_ack_1<= rack(0);
      type_cast_3080_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3080_inst",
        buffer_size => 1,
        in_data_width => 32,
        out_data_width => 32
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => iNsTr_76_2799,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_3080_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3084_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3084_inst_req_0;
      type_cast_3084_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3084_inst_req_1;
      type_cast_3084_inst_ack_1<= rack(0);
      type_cast_3084_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3084_inst",
        buffer_size => 1,
        in_data_width => 32,
        out_data_width => 32
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => xx_xlcssa11_3048,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_3084_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3086_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3086_inst_req_0;
      type_cast_3086_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3086_inst_req_1;
      type_cast_3086_inst_ack_1<= rack(0);
      type_cast_3086_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3086_inst",
        buffer_size => 1,
        in_data_width => 32,
        out_data_width => 32
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tempx_x0x_xphx_xix_xi14_2949,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_3086_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3118_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3118_inst_req_0;
      type_cast_3118_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3118_inst_req_1;
      type_cast_3118_inst_ack_1<= rack(0);
      type_cast_3118_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3118_inst",
        buffer_size => 1,
        in_data_width => 32,
        out_data_width => 32
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => iNsTr_133_3115,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp3x_xix_xi27_3119,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3125_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3125_inst_req_0;
      type_cast_3125_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3125_inst_req_1;
      type_cast_3125_inst_ack_1<= rack(0);
      type_cast_3125_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3125_inst",
        buffer_size => 1,
        in_data_width => 32,
        out_data_width => 32
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp3x_xix_xi27_3119,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_3125_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3144_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3144_inst_req_0;
      type_cast_3144_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3144_inst_req_1;
      type_cast_3144_inst_ack_1<= rack(0);
      type_cast_3144_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3144_inst",
        buffer_size => 1,
        in_data_width => 32,
        out_data_width => 32
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => torque_refx_x0_2190,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp10x_xix_xi_3145,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3148_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3148_inst_req_0;
      type_cast_3148_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3148_inst_req_1;
      type_cast_3148_inst_ack_1<= rack(0);
      type_cast_3148_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3148_inst",
        buffer_size => 1,
        in_data_width => 32,
        out_data_width => 32
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => xx_xop_3141,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => iNsTr_61_3149,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3262_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3262_inst_req_0;
      type_cast_3262_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3262_inst_req_1;
      type_cast_3262_inst_ack_1<= rack(0);
      type_cast_3262_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3262_inst",
        buffer_size => 1,
        in_data_width => 32,
        out_data_width => 32
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => iNsTr_190_3365,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_3262_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3264_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3264_inst_req_0;
      type_cast_3264_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3264_inst_req_1;
      type_cast_3264_inst_ack_1<= rack(0);
      type_cast_3264_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3264_inst",
        buffer_size => 1,
        in_data_width => 32,
        out_data_width => 32
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => iNsTr_94_3211,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_3264_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3268_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3268_inst_req_0;
      type_cast_3268_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3268_inst_req_1;
      type_cast_3268_inst_ack_1<= rack(0);
      type_cast_3268_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3268_inst",
        buffer_size => 1,
        in_data_width => 32,
        out_data_width => 32
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => iNsTr_189_3360,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_3268_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3296_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3296_inst_req_0;
      type_cast_3296_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3296_inst_req_1;
      type_cast_3296_inst_ack_1<= rack(0);
      type_cast_3296_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3296_inst",
        buffer_size => 1,
        in_data_width => 32,
        out_data_width => 32
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => iNsTr_226_3312,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_3296_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3298_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3298_inst_req_0;
      type_cast_3298_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3298_inst_req_1;
      type_cast_3298_inst_ack_1<= rack(0);
      type_cast_3298_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3298_inst",
        buffer_size => 1,
        in_data_width => 32,
        out_data_width => 32
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => iNsTr_97_3229,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_3298_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3302_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3302_inst_req_0;
      type_cast_3302_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3302_inst_req_1;
      type_cast_3302_inst_ack_1<= rack(0);
      type_cast_3302_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3302_inst",
        buffer_size => 1,
        in_data_width => 32,
        out_data_width => 32
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => iNsTr_227_3318,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_3302_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3334_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3334_inst_req_0;
      type_cast_3334_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3334_inst_req_1;
      type_cast_3334_inst_ack_1<= rack(0);
      type_cast_3334_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3334_inst",
        buffer_size => 1,
        in_data_width => 32,
        out_data_width => 32
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => iNsTr_227_3318,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_3334_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3338_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3338_inst_req_0;
      type_cast_3338_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3338_inst_req_1;
      type_cast_3338_inst_ack_1<= rack(0);
      type_cast_3338_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3338_inst",
        buffer_size => 1,
        in_data_width => 32,
        out_data_width => 32
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => iNsTr_226_3312,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_3338_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3345_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3345_inst_req_0;
      type_cast_3345_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3345_inst_req_1;
      type_cast_3345_inst_ack_1<= rack(0);
      type_cast_3345_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3345_inst",
        buffer_size => 1,
        in_data_width => 32,
        out_data_width => 32
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => iNsTr_97_3229,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_3345_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3347_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3347_inst_req_0;
      type_cast_3347_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3347_inst_req_1;
      type_cast_3347_inst_ack_1<= rack(0);
      type_cast_3347_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3347_inst",
        buffer_size => 1,
        in_data_width => 32,
        out_data_width => 32
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => xx_xlcssa7_3335,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_3347_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3354_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3354_inst_req_0;
      type_cast_3354_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3354_inst_req_1;
      type_cast_3354_inst_ack_1<= rack(0);
      type_cast_3354_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3354_inst",
        buffer_size => 1,
        in_data_width => 32,
        out_data_width => 32
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => xx_xlcssa8_3331,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_3354_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3381_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3381_inst_req_0;
      type_cast_3381_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3381_inst_req_1;
      type_cast_3381_inst_ack_1<= rack(0);
      type_cast_3381_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3381_inst",
        buffer_size => 1,
        in_data_width => 32,
        out_data_width => 32
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => iNsTr_189_3360,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_3381_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3391_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3391_inst_req_0;
      type_cast_3391_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3391_inst_req_1;
      type_cast_3391_inst_ack_1<= rack(0);
      type_cast_3391_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3391_inst",
        buffer_size => 1,
        in_data_width => 32,
        out_data_width => 32
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => xx_xlcssa9_3378,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_3391_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3398_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3398_inst_req_0;
      type_cast_3398_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3398_inst_req_1;
      type_cast_3398_inst_ack_1<= rack(0);
      type_cast_3398_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3398_inst",
        buffer_size => 1,
        in_data_width => 32,
        out_data_width => 32
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => xx_x0x_xix_xix_xi_3385,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_3398_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3400_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3400_inst_req_0;
      type_cast_3400_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3400_inst_req_1;
      type_cast_3400_inst_ack_1<= rack(0);
      type_cast_3400_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3400_inst",
        buffer_size => 1,
        in_data_width => 32,
        out_data_width => 32
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => iNsTr_94_3211,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_3400_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3439_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3439_inst_req_0;
      type_cast_3439_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3439_inst_req_1;
      type_cast_3439_inst_ack_1<= rack(0);
      type_cast_3439_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3439_inst",
        buffer_size => 1,
        in_data_width => 32,
        out_data_width => 32
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnextx_xix_xi_3486,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_3439_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3446_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3446_inst_req_0;
      type_cast_3446_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3446_inst_req_1;
      type_cast_3446_inst_ack_1<= rack(0);
      type_cast_3446_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3446_inst",
        buffer_size => 1,
        in_data_width => 32,
        out_data_width => 32
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => iNsTr_194_3455,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_3446_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3448_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3448_inst_req_0;
      type_cast_3448_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3448_inst_req_1;
      type_cast_3448_inst_ack_1<= rack(0);
      type_cast_3448_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3448_inst",
        buffer_size => 1,
        in_data_width => 32,
        out_data_width => 32
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tempx_x0x_xphx_xix_xi_3395,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_3448_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3497_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3497_inst_req_0;
      type_cast_3497_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3497_inst_req_1;
      type_cast_3497_inst_ack_1<= rack(0);
      type_cast_3497_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3497_inst",
        buffer_size => 1,
        in_data_width => 32,
        out_data_width => 32
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => iNsTr_194_3455,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_3497_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3501_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3501_inst_req_0;
      type_cast_3501_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3501_inst_req_1;
      type_cast_3501_inst_ack_1<= rack(0);
      type_cast_3501_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3501_inst",
        buffer_size => 1,
        in_data_width => 32,
        out_data_width => 32
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => iNsTr_193_3436,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_3501_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3524_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3524_inst_req_0;
      type_cast_3524_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3524_inst_req_1;
      type_cast_3524_inst_ack_1<= rack(0);
      type_cast_3524_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3524_inst",
        buffer_size => 1,
        in_data_width => 32,
        out_data_width => 32
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp26x_xix_xi_3518,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_3524_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3526_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3526_inst_req_0;
      type_cast_3526_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3526_inst_req_1;
      type_cast_3526_inst_ack_1<= rack(0);
      type_cast_3526_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3526_inst",
        buffer_size => 1,
        in_data_width => 32,
        out_data_width => 32
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => iNsTr_100_3245,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_3526_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3530_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3530_inst_req_0;
      type_cast_3530_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3530_inst_req_1;
      type_cast_3530_inst_ack_1<= rack(0);
      type_cast_3530_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3530_inst",
        buffer_size => 1,
        in_data_width => 32,
        out_data_width => 32
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => xx_xlcssa6_3494,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_3530_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3532_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3532_inst_req_0;
      type_cast_3532_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3532_inst_req_1;
      type_cast_3532_inst_ack_1<= rack(0);
      type_cast_3532_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3532_inst",
        buffer_size => 1,
        in_data_width => 32,
        out_data_width => 32
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tempx_x0x_xphx_xix_xi_3395,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_3532_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3564_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3564_inst_req_0;
      type_cast_3564_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3564_inst_req_1;
      type_cast_3564_inst_ack_1<= rack(0);
      type_cast_3564_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3564_inst",
        buffer_size => 1,
        in_data_width => 32,
        out_data_width => 32
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => iNsTr_162_3561,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp3x_xix_xi_3565,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3571_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3571_inst_req_0;
      type_cast_3571_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3571_inst_req_1;
      type_cast_3571_inst_ack_1<= rack(0);
      type_cast_3571_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3571_inst",
        buffer_size => 1,
        in_data_width => 32,
        out_data_width => 32
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp3x_xix_xi_3565,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_3571_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3629_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3629_inst_req_0;
      type_cast_3629_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3629_inst_req_1;
      type_cast_3629_inst_ack_1<= rack(0);
      type_cast_3629_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3629_inst",
        buffer_size => 1,
        in_data_width => 32,
        out_data_width => 32
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => iNsTr_85_3597,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_3629_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3690_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3690_inst_req_0;
      type_cast_3690_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3690_inst_req_1;
      type_cast_3690_inst_ack_1<= rack(0);
      type_cast_3690_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3690_inst",
        buffer_size => 1,
        in_data_width => 32,
        out_data_width => 32
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => iNsTr_114_3647,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_3690_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3700_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3700_inst_req_0;
      type_cast_3700_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3700_inst_req_1;
      type_cast_3700_inst_ack_1<= rack(0);
      type_cast_3700_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3700_inst",
        buffer_size => 1,
        in_data_width => 32,
        out_data_width => 32
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp10x_xi55x_xin_3687,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp10x_xi55_3701,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3725_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3725_inst_req_0;
      type_cast_3725_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3725_inst_req_1;
      type_cast_3725_inst_ack_1<= rack(0);
      type_cast_3725_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3725_inst",
        buffer_size => 1,
        in_data_width => 32,
        out_data_width => 32
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => iNsTr_213_3831,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_3725_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3727_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3727_inst_req_0;
      type_cast_3727_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3727_inst_req_1;
      type_cast_3727_inst_ack_1<= rack(0);
      type_cast_3727_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3727_inst",
        buffer_size => 1,
        in_data_width => 32,
        out_data_width => 32
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => iNsTr_149_3719,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_3727_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3731_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3731_inst_req_0;
      type_cast_3731_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3731_inst_req_1;
      type_cast_3731_inst_ack_1<= rack(0);
      type_cast_3731_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3731_inst",
        buffer_size => 1,
        in_data_width => 32,
        out_data_width => 32
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => iNsTr_212_3826,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_3731_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3760_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3760_inst_req_0;
      type_cast_3760_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3760_inst_req_1;
      type_cast_3760_inst_ack_1<= rack(0);
      type_cast_3760_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3760_inst",
        buffer_size => 1,
        in_data_width => 32,
        out_data_width => 32
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => iNsTr_234_3777,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_3760_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3767_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3767_inst_req_0;
      type_cast_3767_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3767_inst_req_1;
      type_cast_3767_inst_ack_1<= rack(0);
      type_cast_3767_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3767_inst",
        buffer_size => 1,
        in_data_width => 32,
        out_data_width => 32
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => iNsTr_235_3783,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_3767_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3799_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3799_inst_req_0;
      type_cast_3799_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3799_inst_req_1;
      type_cast_3799_inst_ack_1<= rack(0);
      type_cast_3799_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3799_inst",
        buffer_size => 1,
        in_data_width => 32,
        out_data_width => 32
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => iNsTr_235_3783,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_3799_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3803_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3803_inst_req_0;
      type_cast_3803_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3803_inst_req_1;
      type_cast_3803_inst_ack_1<= rack(0);
      type_cast_3803_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3803_inst",
        buffer_size => 1,
        in_data_width => 32,
        out_data_width => 32
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => iNsTr_234_3777,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_3803_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3813_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3813_inst_req_0;
      type_cast_3813_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3813_inst_req_1;
      type_cast_3813_inst_ack_1<= rack(0);
      type_cast_3813_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3813_inst",
        buffer_size => 1,
        in_data_width => 32,
        out_data_width => 32
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => xx_xlcssa2_3800,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_3813_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3820_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3820_inst_req_0;
      type_cast_3820_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3820_inst_req_1;
      type_cast_3820_inst_ack_1<= rack(0);
      type_cast_3820_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3820_inst",
        buffer_size => 1,
        in_data_width => 32,
        out_data_width => 32
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => xx_xlcssa3_3796,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_3820_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3848_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3848_inst_req_0;
      type_cast_3848_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3848_inst_req_1;
      type_cast_3848_inst_ack_1<= rack(0);
      type_cast_3848_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3848_inst",
        buffer_size => 1,
        in_data_width => 32,
        out_data_width => 32
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => iNsTr_212_3826,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_3848_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3911_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3911_inst_req_0;
      type_cast_3911_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3911_inst_req_1;
      type_cast_3911_inst_ack_1<= rack(0);
      type_cast_3911_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3911_inst",
        buffer_size => 1,
        in_data_width => 32,
        out_data_width => 32
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnextx_xi_3958,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_3911_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3918_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3918_inst_req_0;
      type_cast_3918_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3918_inst_req_1;
      type_cast_3918_inst_ack_1<= rack(0);
      type_cast_3918_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3918_inst",
        buffer_size => 1,
        in_data_width => 32,
        out_data_width => 32
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => iNsTr_256_3927,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_3918_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3920_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3920_inst_req_0;
      type_cast_3920_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3920_inst_req_1;
      type_cast_3920_inst_ack_1<= rack(0);
      type_cast_3920_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3920_inst",
        buffer_size => 1,
        in_data_width => 32,
        out_data_width => 32
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => xx_xlcssa4_3845,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_3920_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3969_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3969_inst_req_0;
      type_cast_3969_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3969_inst_req_1;
      type_cast_3969_inst_ack_1<= rack(0);
      type_cast_3969_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3969_inst",
        buffer_size => 1,
        in_data_width => 32,
        out_data_width => 32
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => iNsTr_256_3927,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_3969_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3973_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3973_inst_req_0;
      type_cast_3973_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3973_inst_req_1;
      type_cast_3973_inst_ack_1<= rack(0);
      type_cast_3973_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3973_inst",
        buffer_size => 1,
        in_data_width => 32,
        out_data_width => 32
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => iNsTr_255_3908,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_3973_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3991_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3991_inst_req_0;
      type_cast_3991_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3991_inst_req_1;
      type_cast_3991_inst_ack_1<= rack(0);
      type_cast_3991_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3991_inst",
        buffer_size => 1,
        in_data_width => 32,
        out_data_width => 32
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp26x_xi_3985,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_3991_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3993_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3993_inst_req_0;
      type_cast_3993_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3993_inst_req_1;
      type_cast_3993_inst_ack_1<= rack(0);
      type_cast_3993_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3993_inst",
        buffer_size => 1,
        in_data_width => 32,
        out_data_width => 32
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => iNsTr_241_3873,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_3993_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3997_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3997_inst_req_0;
      type_cast_3997_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3997_inst_req_1;
      type_cast_3997_inst_ack_1<= rack(0);
      type_cast_3997_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3997_inst",
        buffer_size => 1,
        in_data_width => 32,
        out_data_width => 32
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => xx_xlcssa1_3966,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_3997_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3999_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3999_inst_req_0;
      type_cast_3999_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3999_inst_req_1;
      type_cast_3999_inst_ack_1<= rack(0);
      type_cast_3999_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3999_inst",
        buffer_size => 1,
        in_data_width => 32,
        out_data_width => 32
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => xx_xlcssa4_3845,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_3999_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_4031_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_4031_inst_req_0;
      type_cast_4031_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_4031_inst_req_1;
      type_cast_4031_inst_ack_1<= rack(0);
      type_cast_4031_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_4031_inst",
        buffer_size => 1,
        in_data_width => 32,
        out_data_width => 32
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => iNsTr_253_4028,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp3x_xi_4032,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_4038_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_4038_inst_req_0;
      type_cast_4038_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_4038_inst_req_1;
      type_cast_4038_inst_ack_1<= rack(0);
      type_cast_4038_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_4038_inst",
        buffer_size => 1,
        in_data_width => 32,
        out_data_width => 32
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp3x_xi_4032,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_4038_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    if_stmt_2112_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= iNsTr_14_2111;
      branch_instance: BranchBase -- 
        generic map( condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2112_branch_req_0,
          ack0 => if_stmt_2112_branch_ack_0,
          ack1 => if_stmt_2112_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_2125_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= iNsTr_20_2124;
      branch_instance: BranchBase -- 
        generic map( condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2125_branch_req_0,
          ack0 => if_stmt_2125_branch_ack_0,
          ack1 => if_stmt_2125_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_2162_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= iNsTr_18_2161;
      branch_instance: BranchBase -- 
        generic map( condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2162_branch_req_0,
          ack0 => if_stmt_2162_branch_ack_0,
          ack1 => if_stmt_2162_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_2175_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= iNsTr_25_2174;
      branch_instance: BranchBase -- 
        generic map( condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2175_branch_req_0,
          ack0 => if_stmt_2175_branch_ack_0,
          ack1 => if_stmt_2175_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_2211_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= iNsTr_23_2210;
      branch_instance: BranchBase -- 
        generic map( condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2211_branch_req_0,
          ack0 => if_stmt_2211_branch_ack_0,
          ack1 => if_stmt_2211_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_2224_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= iNsTr_28_2223;
      branch_instance: BranchBase -- 
        generic map( condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2224_branch_req_0,
          ack0 => if_stmt_2224_branch_ack_0,
          ack1 => if_stmt_2224_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_2257_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= iNsTr_36_2256;
      branch_instance: BranchBase -- 
        generic map( condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2257_branch_req_0,
          ack0 => if_stmt_2257_branch_ack_0,
          ack1 => if_stmt_2257_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_2343_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= iNsTr_33_2342;
      branch_instance: BranchBase -- 
        generic map( condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2343_branch_req_0,
          ack0 => if_stmt_2343_branch_ack_0,
          ack1 => if_stmt_2343_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_2396_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= iNsTr_79_2395;
      branch_instance: BranchBase -- 
        generic map( condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2396_branch_req_0,
          ack0 => if_stmt_2396_branch_ack_0,
          ack1 => if_stmt_2396_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_2437_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= iNsTr_137_2436;
      branch_instance: BranchBase -- 
        generic map( condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2437_branch_req_0,
          ack0 => if_stmt_2437_branch_ack_0,
          ack1 => if_stmt_2437_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_2486_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= iNsTr_111_2485;
      branch_instance: BranchBase -- 
        generic map( condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2486_branch_req_0,
          ack0 => if_stmt_2486_branch_ack_0,
          ack1 => if_stmt_2486_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_2547_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= orx_xcond11x_xix_xi40_2546;
      branch_instance: BranchBase -- 
        generic map( condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2547_branch_req_0,
          ack0 => if_stmt_2547_branch_ack_0,
          ack1 => if_stmt_2547_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_2607_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= orx_xcondx_xix_xi43_2600;
      branch_instance: BranchBase -- 
        generic map( condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2607_branch_req_0,
          ack0 => if_stmt_2607_branch_ack_0,
          ack1 => if_stmt_2607_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_2717_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= iNsTr_45_2716;
      branch_instance: BranchBase -- 
        generic map( condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2717_branch_req_0,
          ack0 => if_stmt_2717_branch_ack_0,
          ack1 => if_stmt_2717_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_2838_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= iNsTr_126_2837;
      branch_instance: BranchBase -- 
        generic map( condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2838_branch_req_0,
          ack0 => if_stmt_2838_branch_ack_0,
          ack1 => if_stmt_2838_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_2878_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= iNsTr_201_2877;
      branch_instance: BranchBase -- 
        generic map( condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2878_branch_req_0,
          ack0 => if_stmt_2878_branch_ack_0,
          ack1 => if_stmt_2878_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_2925_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= iNsTr_167_2924;
      branch_instance: BranchBase -- 
        generic map( condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2925_branch_req_0,
          ack0 => if_stmt_2925_branch_ack_0,
          ack1 => if_stmt_2925_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_2981_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= orx_xcond11x_xix_xi15_2980;
      branch_instance: BranchBase -- 
        generic map( condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2981_branch_req_0,
          ack0 => if_stmt_2981_branch_ack_0,
          ack1 => if_stmt_2981_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_3041_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= orx_xcondx_xix_xi18_3034;
      branch_instance: BranchBase -- 
        generic map( condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_3041_branch_req_0,
          ack0 => if_stmt_3041_branch_ack_0,
          ack1 => if_stmt_3041_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_3163_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= iNsTr_62_3162;
      branch_instance: BranchBase -- 
        generic map( condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_3163_branch_req_0,
          ack0 => if_stmt_3163_branch_ack_0,
          ack1 => if_stmt_3163_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_3284_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= iNsTr_155_3283;
      branch_instance: BranchBase -- 
        generic map( condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_3284_branch_req_0,
          ack0 => if_stmt_3284_branch_ack_0,
          ack1 => if_stmt_3284_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_3324_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= iNsTr_228_3323;
      branch_instance: BranchBase -- 
        generic map( condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_3324_branch_req_0,
          ack0 => if_stmt_3324_branch_ack_0,
          ack1 => if_stmt_3324_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_3371_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= iNsTr_191_3370;
      branch_instance: BranchBase -- 
        generic map( condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_3371_branch_req_0,
          ack0 => if_stmt_3371_branch_ack_0,
          ack1 => if_stmt_3371_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_3427_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= orx_xcond11x_xix_xi_3426;
      branch_instance: BranchBase -- 
        generic map( condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_3427_branch_req_0,
          ack0 => if_stmt_3427_branch_ack_0,
          ack1 => if_stmt_3427_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_3487_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= orx_xcondx_xix_xi_3480;
      branch_instance: BranchBase -- 
        generic map( condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_3487_branch_req_0,
          ack0 => if_stmt_3487_branch_ack_0,
          ack1 => if_stmt_3487_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_3604_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= iNsTr_86_3603;
      branch_instance: BranchBase -- 
        generic map( condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_3604_branch_req_0,
          ack0 => if_stmt_3604_branch_ack_0,
          ack1 => if_stmt_3604_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_3617_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= iNsTr_117_3616;
      branch_instance: BranchBase -- 
        generic map( condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_3617_branch_req_0,
          ack0 => if_stmt_3617_branch_ack_0,
          ack1 => if_stmt_3617_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_3654_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= iNsTr_115_3653;
      branch_instance: BranchBase -- 
        generic map( condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_3654_branch_req_0,
          ack0 => if_stmt_3654_branch_ack_0,
          ack1 => if_stmt_3654_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_3667_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= iNsTr_151_3666;
      branch_instance: BranchBase -- 
        generic map( condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_3667_branch_req_0,
          ack0 => if_stmt_3667_branch_ack_0,
          ack1 => if_stmt_3667_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_3680_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= iNsTr_186_3679;
      branch_instance: BranchBase -- 
        generic map( condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_3680_branch_req_0,
          ack0 => if_stmt_3680_branch_ack_0,
          ack1 => if_stmt_3680_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_3748_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= iNsTr_184_3747;
      branch_instance: BranchBase -- 
        generic map( condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_3748_branch_req_0,
          ack0 => if_stmt_3748_branch_ack_0,
          ack1 => if_stmt_3748_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_3789_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= iNsTr_236_3788;
      branch_instance: BranchBase -- 
        generic map( condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_3789_branch_req_0,
          ack0 => if_stmt_3789_branch_ack_0,
          ack1 => if_stmt_3789_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_3838_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= iNsTr_214_3837;
      branch_instance: BranchBase -- 
        generic map( condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_3838_branch_req_0,
          ack0 => if_stmt_3838_branch_ack_0,
          ack1 => if_stmt_3838_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_3899_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= orx_xcond11x_xi_3898;
      branch_instance: BranchBase -- 
        generic map( condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_3899_branch_req_0,
          ack0 => if_stmt_3899_branch_ack_0,
          ack1 => if_stmt_3899_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_3959_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= orx_xcondx_xi_3952;
      branch_instance: BranchBase -- 
        generic map( condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_3959_branch_req_0,
          ack0 => if_stmt_3959_branch_ack_0,
          ack1 => if_stmt_3959_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    switch_stmt_2800_branch_0: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= expr_2802_wire_constant_cmp;
      branch_instance: BranchBase -- 
        generic map( condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => switch_stmt_2800_branch_0_req_0,
          ack0 => open,
          ack1 => switch_stmt_2800_branch_0_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    switch_stmt_2800_branch_1: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= expr_2805_wire_constant_cmp;
      branch_instance: BranchBase -- 
        generic map( condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => switch_stmt_2800_branch_1_req_0,
          ack0 => open,
          ack1 => switch_stmt_2800_branch_1_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    switch_stmt_2800_branch_default: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(1 downto 0);
      begin 
      condition_sig <= expr_2802_wire_constant_cmp & expr_2805_wire_constant_cmp;
      branch_instance: BranchBase -- 
        generic map( condition_width => 2)
        port map( -- 
          condition => condition_sig,
          req => switch_stmt_2800_branch_default_req_0,
          ack0 => switch_stmt_2800_branch_default_ack_0,
          ack1 => open,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    switch_stmt_3246_branch_0: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= expr_3248_wire_constant_cmp;
      branch_instance: BranchBase -- 
        generic map( condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => switch_stmt_3246_branch_0_req_0,
          ack0 => open,
          ack1 => switch_stmt_3246_branch_0_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    switch_stmt_3246_branch_1: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= expr_3251_wire_constant_cmp;
      branch_instance: BranchBase -- 
        generic map( condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => switch_stmt_3246_branch_1_req_0,
          ack0 => open,
          ack1 => switch_stmt_3246_branch_1_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    switch_stmt_3246_branch_default: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(1 downto 0);
      begin 
      condition_sig <= expr_3248_wire_constant_cmp & expr_3251_wire_constant_cmp;
      branch_instance: BranchBase -- 
        generic map( condition_width => 2)
        port map( -- 
          condition => condition_sig,
          req => switch_stmt_3246_branch_default_req_0,
          ack0 => switch_stmt_3246_branch_default_ack_0,
          ack1 => open,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- shared split operator group (0) : ADD_f32_f32_2093_inst ADD_f32_f32_2241_inst ADD_f32_f32_2154_inst ADD_f32_f32_2274_inst ADD_f32_f32_2331_inst ADD_f32_f32_2294_inst ADD_f32_f32_3590_inst ADD_f32_f32_3646_inst 
    ApFloatAdd_group_0: Block -- 
      signal data_in: std_logic_vector(511 downto 0);
      signal data_out: std_logic_vector(255 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 7 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 7 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 7 downto 0);
      signal guard_vector : std_logic_vector( 7 downto 0);
      constant inBUFs : IntegerArray(7 downto 0) := (7 => 1, 6 => 1, 5 => 1, 4 => 1, 3 => 1, 2 => 1, 1 => 1, 0 => 1);
      constant outBUFs : IntegerArray(7 downto 0) := (7 => 1, 6 => 1, 5 => 1, 4 => 1, 3 => 1, 2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(7 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false);
      constant guardBuffering: IntegerArray(7 downto 0)  := (0 => 1, 1 => 1, 2 => 1, 3 => 1, 4 => 1, 5 => 1, 6 => 1, 7 => 1);
      -- 
    begin -- 
      data_in <= iNsTr_10_2089 & int_speed_errx_x0_2059 & iNsTr_38_2236 & type_cast_2240_wire_constant & int_speed_errx_x1_2134 & iNsTr_16_2150 & iNsTr_55_2269 & type_cast_2273_wire_constant & iNsTr_31_2327 & iNsTr_30_2321 & iNsTr_51_2289 & type_cast_2293_wire_constant & iNsTr_83_3586 & int_flux_errx_x0_2052 & int_flux_errx_x1_3626 & iNsTr_113_3642;
      iNsTr_11_2094 <= data_out(255 downto 224);
      iNsTr_39_2242 <= data_out(223 downto 192);
      iNsTr_17_2155 <= data_out(191 downto 160);
      iNsTr_56_2275 <= data_out(159 downto 128);
      iNsTr_32_2332 <= data_out(127 downto 96);
      iNsTr_52_2295 <= data_out(95 downto 64);
      iNsTr_84_3591 <= data_out(63 downto 32);
      iNsTr_114_3647 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      reqL_unguarded(7) <= ADD_f32_f32_2093_inst_req_0;
      reqL_unguarded(6) <= ADD_f32_f32_2241_inst_req_0;
      reqL_unguarded(5) <= ADD_f32_f32_2154_inst_req_0;
      reqL_unguarded(4) <= ADD_f32_f32_2274_inst_req_0;
      reqL_unguarded(3) <= ADD_f32_f32_2331_inst_req_0;
      reqL_unguarded(2) <= ADD_f32_f32_2294_inst_req_0;
      reqL_unguarded(1) <= ADD_f32_f32_3590_inst_req_0;
      reqL_unguarded(0) <= ADD_f32_f32_3646_inst_req_0;
      ADD_f32_f32_2093_inst_ack_0 <= ackL_unguarded(7);
      ADD_f32_f32_2241_inst_ack_0 <= ackL_unguarded(6);
      ADD_f32_f32_2154_inst_ack_0 <= ackL_unguarded(5);
      ADD_f32_f32_2274_inst_ack_0 <= ackL_unguarded(4);
      ADD_f32_f32_2331_inst_ack_0 <= ackL_unguarded(3);
      ADD_f32_f32_2294_inst_ack_0 <= ackL_unguarded(2);
      ADD_f32_f32_3590_inst_ack_0 <= ackL_unguarded(1);
      ADD_f32_f32_3646_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(7) <= ADD_f32_f32_2093_inst_req_1;
      reqR_unguarded(6) <= ADD_f32_f32_2241_inst_req_1;
      reqR_unguarded(5) <= ADD_f32_f32_2154_inst_req_1;
      reqR_unguarded(4) <= ADD_f32_f32_2274_inst_req_1;
      reqR_unguarded(3) <= ADD_f32_f32_2331_inst_req_1;
      reqR_unguarded(2) <= ADD_f32_f32_2294_inst_req_1;
      reqR_unguarded(1) <= ADD_f32_f32_3590_inst_req_1;
      reqR_unguarded(0) <= ADD_f32_f32_3646_inst_req_1;
      ADD_f32_f32_2093_inst_ack_1 <= ackR_unguarded(7);
      ADD_f32_f32_2241_inst_ack_1 <= ackR_unguarded(6);
      ADD_f32_f32_2154_inst_ack_1 <= ackR_unguarded(5);
      ADD_f32_f32_2274_inst_ack_1 <= ackR_unguarded(4);
      ADD_f32_f32_2331_inst_ack_1 <= ackR_unguarded(3);
      ADD_f32_f32_2294_inst_ack_1 <= ackR_unguarded(2);
      ADD_f32_f32_3590_inst_ack_1 <= ackR_unguarded(1);
      ADD_f32_f32_3646_inst_ack_1 <= ackR_unguarded(0);
      ApFloatAdd_group_0_accessRegulator_0: access_regulator_base generic map (name => "ApFloatAdd_group_0_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      ApFloatAdd_group_0_accessRegulator_1: access_regulator_base generic map (name => "ApFloatAdd_group_0_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      ApFloatAdd_group_0_accessRegulator_2: access_regulator_base generic map (name => "ApFloatAdd_group_0_accessRegulator_2", num_slots => 1) -- 
        port map (req => reqL_unregulated(2), -- 
          ack => ackL_unregulated(2),
          regulated_req => reqL(2),
          regulated_ack => ackL(2),
          release_req => reqR(2),
          release_ack => ackR(2),
          clk => clk, reset => reset); -- 
      ApFloatAdd_group_0_accessRegulator_3: access_regulator_base generic map (name => "ApFloatAdd_group_0_accessRegulator_3", num_slots => 1) -- 
        port map (req => reqL_unregulated(3), -- 
          ack => ackL_unregulated(3),
          regulated_req => reqL(3),
          regulated_ack => ackL(3),
          release_req => reqR(3),
          release_ack => ackR(3),
          clk => clk, reset => reset); -- 
      ApFloatAdd_group_0_accessRegulator_4: access_regulator_base generic map (name => "ApFloatAdd_group_0_accessRegulator_4", num_slots => 1) -- 
        port map (req => reqL_unregulated(4), -- 
          ack => ackL_unregulated(4),
          regulated_req => reqL(4),
          regulated_ack => ackL(4),
          release_req => reqR(4),
          release_ack => ackR(4),
          clk => clk, reset => reset); -- 
      ApFloatAdd_group_0_accessRegulator_5: access_regulator_base generic map (name => "ApFloatAdd_group_0_accessRegulator_5", num_slots => 1) -- 
        port map (req => reqL_unregulated(5), -- 
          ack => ackL_unregulated(5),
          regulated_req => reqL(5),
          regulated_ack => ackL(5),
          release_req => reqR(5),
          release_ack => ackR(5),
          clk => clk, reset => reset); -- 
      ApFloatAdd_group_0_accessRegulator_6: access_regulator_base generic map (name => "ApFloatAdd_group_0_accessRegulator_6", num_slots => 1) -- 
        port map (req => reqL_unregulated(6), -- 
          ack => ackL_unregulated(6),
          regulated_req => reqL(6),
          regulated_ack => ackL(6),
          release_req => reqR(6),
          release_ack => ackR(6),
          clk => clk, reset => reset); -- 
      ApFloatAdd_group_0_accessRegulator_7: access_regulator_base generic map (name => "ApFloatAdd_group_0_accessRegulator_7", num_slots => 1) -- 
        port map (req => reqL_unregulated(7), -- 
          ack => ackL_unregulated(7),
          regulated_req => reqL(7),
          regulated_ack => ackL(7),
          release_req => reqR(7),
          release_ack => ackR(7),
          clk => clk, reset => reset); -- 
      gI: SplitGuardInterface generic map(nreqs => 8, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      PipedFpOp: PipelinedFPOperator -- 
        generic map( -- 
          name => "ApFloatAdd_group_0",
          operator_id => "ApFloatAdd",
          exponent_width => 8,
          fraction_width => 23, 
          no_arbitration => false,
          num_reqs => 8,
          use_input_buffering => true,
          detailed_buffering_per_input => inBUFs,
          detailed_buffering_per_output => outBUFs -- 
        )
        port map ( reqL => reqL , ackL => ackL, reqR => reqR, ackR => ackR, dataL => data_in, dataR => data_out, clk => clk, reset => reset); -- 
      -- 
    end Block; -- split operator group 0
    -- shared split operator group (1) : ADD_u32_u32_2473_inst 
    ApIntAdd_group_1: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= curr_quotientx_x0x_xlcssax_xix_xix_xi38_2462 & quotientx_x05x_xix_xix_xi32_2376;
      iNsTr_109_2474 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ADD_u32_u32_2473_inst_req_0;
      ADD_u32_u32_2473_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ADD_u32_u32_2473_inst_req_1;
      ADD_u32_u32_2473_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_1",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 1
    -- shared split operator group (2) : ADD_u32_u32_2520_inst 
    ApIntAdd_group_2: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= iNsTr_141_2515;
      iNsTr_142_2521 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ADD_u32_u32_2520_inst_req_0;
      ADD_u32_u32_2520_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ADD_u32_u32_2520_inst_req_1;
      ADD_u32_u32_2520_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_2",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "11111111111111111111111101111011",
          constant_width => 32,
          buffering  => 1,
          flow_through => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 2
    -- shared split operator group (3) : ADD_u32_u32_2605_inst 
    ApIntAdd_group_3: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= iNsTr_205_2556;
      indvarx_xnextx_xix_xi44_2606 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ADD_u32_u32_2605_inst_req_0;
      ADD_u32_u32_2605_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ADD_u32_u32_2605_inst_req_1;
      ADD_u32_u32_2605_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_3",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000001",
          constant_width => 32,
          buffering  => 1,
          flow_through => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 3
    -- shared split operator group (4) : ADD_u32_u32_2627_inst 
    ApIntAdd_group_4: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= iNsTr_141_2515;
      tmp25x_xix_xi46_2628 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ADD_u32_u32_2627_inst_req_0;
      ADD_u32_u32_2627_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ADD_u32_u32_2627_inst_req_1;
      ADD_u32_u32_2627_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_4",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "11111111111111111111111101111010",
          constant_width => 32,
          buffering  => 1,
          flow_through => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 4
    -- shared split operator group (5) : ADD_u32_u32_2665_inst 
    ApIntAdd_group_5: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= iNsTr_178_2660;
      iNsTr_179_2666 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ADD_u32_u32_2665_inst_req_0;
      ADD_u32_u32_2665_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ADD_u32_u32_2665_inst_req_1;
      ADD_u32_u32_2665_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_5",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "01000100000000000000000000000000",
          constant_width => 32,
          buffering  => 1,
          flow_through => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 5
    -- shared split operator group (6) : ADD_u32_u32_2913_inst 
    ApIntAdd_group_6: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= curr_quotientx_x0x_xlcssax_xix_xix_xi10_2902 & quotientx_x05x_xix_xix_xi4_2819;
      iNsTr_165_2914 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ADD_u32_u32_2913_inst_req_0;
      ADD_u32_u32_2913_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ADD_u32_u32_2913_inst_req_1;
      ADD_u32_u32_2913_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_6",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 6
    -- shared split operator group (7) : ADD_u32_u32_3039_inst 
    ApIntAdd_group_7: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= iNsTr_169_2990;
      indvarx_xnextx_xix_xi19_3040 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ADD_u32_u32_3039_inst_req_0;
      ADD_u32_u32_3039_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ADD_u32_u32_3039_inst_req_1;
      ADD_u32_u32_3039_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_7",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000001",
          constant_width => 32,
          buffering  => 1,
          flow_through => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 7
    -- shared split operator group (8) : ADD_u32_u32_3061_inst 
    ApIntAdd_group_8: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= iNsTr_65_2735;
      tmp21x_xix_xi21_3062 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ADD_u32_u32_3061_inst_req_0;
      ADD_u32_u32_3061_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ADD_u32_u32_3061_inst_req_1;
      ADD_u32_u32_3061_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_8",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "11111111111111111111111111111111",
          constant_width => 32,
          buffering  => 1,
          flow_through => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 8
    -- shared split operator group (9) : ADD_u32_u32_3104_inst 
    ApIntAdd_group_9: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= iNsTr_130_3099;
      iNsTr_131_3105 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ADD_u32_u32_3104_inst_req_0;
      ADD_u32_u32_3104_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ADD_u32_u32_3104_inst_req_1;
      ADD_u32_u32_3104_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_9",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "01000100000000000000000000000000",
          constant_width => 32,
          buffering  => 1,
          flow_through => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 9
    -- shared split operator group (10) : ADD_u32_u32_3359_inst 
    ApIntAdd_group_10: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= curr_quotientx_x0x_xlcssax_xix_xix_xi_3348 & quotientx_x05x_xix_xix_xi_3265;
      iNsTr_189_3360 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ADD_u32_u32_3359_inst_req_0;
      ADD_u32_u32_3359_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ADD_u32_u32_3359_inst_req_1;
      ADD_u32_u32_3359_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_10",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 10
    -- shared split operator group (11) : ADD_u32_u32_3485_inst 
    ApIntAdd_group_11: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= iNsTr_193_3436;
      indvarx_xnextx_xix_xi_3486 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ADD_u32_u32_3485_inst_req_0;
      ADD_u32_u32_3485_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ADD_u32_u32_3485_inst_req_1;
      ADD_u32_u32_3485_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_11",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000001",
          constant_width => 32,
          buffering  => 1,
          flow_through => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 11
    -- shared split operator group (12) : ADD_u32_u32_3507_inst 
    ApIntAdd_group_12: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= iNsTr_89_3181;
      tmp21x_xix_xi_3508 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ADD_u32_u32_3507_inst_req_0;
      ADD_u32_u32_3507_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ADD_u32_u32_3507_inst_req_1;
      ADD_u32_u32_3507_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_12",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "11111111111111111111111111111111",
          constant_width => 32,
          buffering  => 1,
          flow_through => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 12
    -- shared split operator group (13) : ADD_u32_u32_3550_inst 
    ApIntAdd_group_13: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= iNsTr_159_3545;
      iNsTr_160_3551 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ADD_u32_u32_3550_inst_req_0;
      ADD_u32_u32_3550_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ADD_u32_u32_3550_inst_req_1;
      ADD_u32_u32_3550_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_13",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "01000100000000000000000000000000",
          constant_width => 32,
          buffering  => 1,
          flow_through => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 13
    -- shared split operator group (14) : ADD_u32_u32_3825_inst 
    ApIntAdd_group_14: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= curr_quotientx_x0x_xlcssax_xix_xi_3814 & quotientx_x05x_xix_xi_3728;
      iNsTr_212_3826 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ADD_u32_u32_3825_inst_req_0;
      ADD_u32_u32_3825_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ADD_u32_u32_3825_inst_req_1;
      ADD_u32_u32_3825_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_14",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 14
    -- shared split operator group (15) : ADD_u32_u32_3872_inst 
    ApIntAdd_group_15: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= iNsTr_240_3867;
      iNsTr_241_3873 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ADD_u32_u32_3872_inst_req_0;
      ADD_u32_u32_3872_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ADD_u32_u32_3872_inst_req_1;
      ADD_u32_u32_3872_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_15",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "11111111111111111111111101111011",
          constant_width => 32,
          buffering  => 1,
          flow_through => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 15
    -- shared split operator group (16) : ADD_u32_u32_3957_inst 
    ApIntAdd_group_16: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= iNsTr_255_3908;
      indvarx_xnextx_xi_3958 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ADD_u32_u32_3957_inst_req_0;
      ADD_u32_u32_3957_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ADD_u32_u32_3957_inst_req_1;
      ADD_u32_u32_3957_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_16",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000001",
          constant_width => 32,
          buffering  => 1,
          flow_through => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 16
    -- shared split operator group (17) : ADD_u32_u32_3979_inst 
    ApIntAdd_group_17: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= iNsTr_240_3867;
      tmp25x_xi_3980 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ADD_u32_u32_3979_inst_req_0;
      ADD_u32_u32_3979_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ADD_u32_u32_3979_inst_req_1;
      ADD_u32_u32_3979_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_17",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "11111111111111111111111101111010",
          constant_width => 32,
          buffering  => 1,
          flow_through => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 17
    -- shared split operator group (18) : ADD_u32_u32_4017_inst 
    ApIntAdd_group_18: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= iNsTr_250_4012;
      iNsTr_251_4018 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ADD_u32_u32_4017_inst_req_0;
      ADD_u32_u32_4017_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ADD_u32_u32_4017_inst_req_1;
      ADD_u32_u32_4017_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_18",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "01000100000000000000000000000000",
          constant_width => 32,
          buffering  => 1,
          flow_through => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 18
    -- shared split operator group (19) : AND_u1_u1_2545_inst 
    ApIntAnd_group_19: Block -- 
      signal data_in: std_logic_vector(1 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= iNsTr_144_2533 & iNsTr_145_2541;
      orx_xcond11x_xix_xi40_2546 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= AND_u1_u1_2545_inst_req_0;
      AND_u1_u1_2545_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= AND_u1_u1_2545_inst_req_1;
      AND_u1_u1_2545_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAnd",
          name => "ApIntAnd_group_19",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 1,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 1, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 19
    -- shared split operator group (20) : AND_u1_u1_2599_inst 
    ApIntAnd_group_20: Block -- 
      signal data_in: std_logic_vector(1 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= iNsTr_208_2587 & iNsTr_209_2595;
      orx_xcondx_xix_xi43_2600 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= AND_u1_u1_2599_inst_req_0;
      AND_u1_u1_2599_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= AND_u1_u1_2599_inst_req_1;
      AND_u1_u1_2599_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAnd",
          name => "ApIntAnd_group_20",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 1,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 1, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 20
    -- shared split operator group (21) : AND_u1_u1_2979_inst 
    ApIntAnd_group_21: Block -- 
      signal data_in: std_logic_vector(1 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= iNsTr_105_2967 & iNsTr_106_2975;
      orx_xcond11x_xix_xi15_2980 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= AND_u1_u1_2979_inst_req_0;
      AND_u1_u1_2979_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= AND_u1_u1_2979_inst_req_1;
      AND_u1_u1_2979_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAnd",
          name => "ApIntAnd_group_21",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 1,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 1, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 21
    -- shared split operator group (22) : AND_u1_u1_3033_inst 
    ApIntAnd_group_22: Block -- 
      signal data_in: std_logic_vector(1 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= iNsTr_172_3021 & iNsTr_173_3029;
      orx_xcondx_xix_xi18_3034 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= AND_u1_u1_3033_inst_req_0;
      AND_u1_u1_3033_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= AND_u1_u1_3033_inst_req_1;
      AND_u1_u1_3033_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAnd",
          name => "ApIntAnd_group_22",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 1,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 1, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 22
    -- shared split operator group (23) : AND_u1_u1_3425_inst 
    ApIntAnd_group_23: Block -- 
      signal data_in: std_logic_vector(1 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= iNsTr_122_3413 & iNsTr_123_3421;
      orx_xcond11x_xix_xi_3426 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= AND_u1_u1_3425_inst_req_0;
      AND_u1_u1_3425_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= AND_u1_u1_3425_inst_req_1;
      AND_u1_u1_3425_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAnd",
          name => "ApIntAnd_group_23",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 1,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 1, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 23
    -- shared split operator group (24) : AND_u1_u1_3479_inst 
    ApIntAnd_group_24: Block -- 
      signal data_in: std_logic_vector(1 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= iNsTr_196_3467 & iNsTr_197_3475;
      orx_xcondx_xix_xi_3480 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= AND_u1_u1_3479_inst_req_0;
      AND_u1_u1_3479_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= AND_u1_u1_3479_inst_req_1;
      AND_u1_u1_3479_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAnd",
          name => "ApIntAnd_group_24",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 1,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 1, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 24
    -- shared split operator group (25) : AND_u1_u1_3897_inst 
    ApIntAnd_group_25: Block -- 
      signal data_in: std_logic_vector(1 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= iNsTr_243_3885 & iNsTr_244_3893;
      orx_xcond11x_xi_3898 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= AND_u1_u1_3897_inst_req_0;
      AND_u1_u1_3897_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= AND_u1_u1_3897_inst_req_1;
      AND_u1_u1_3897_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAnd",
          name => "ApIntAnd_group_25",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 1,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 1, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 25
    -- shared split operator group (26) : AND_u1_u1_3951_inst 
    ApIntAnd_group_26: Block -- 
      signal data_in: std_logic_vector(1 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= iNsTr_258_3939 & iNsTr_259_3947;
      orx_xcondx_xi_3952 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= AND_u1_u1_3951_inst_req_0;
      AND_u1_u1_3951_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= AND_u1_u1_3951_inst_req_1;
      AND_u1_u1_3951_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAnd",
          name => "ApIntAnd_group_26",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 1,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 1, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 26
    -- shared split operator group (27) : AND_u32_u32_2360_inst 
    ApIntAnd_group_27: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= iNsTr_47_2355;
      iNsTr_48_2361 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= AND_u32_u32_2360_inst_req_0;
      AND_u32_u32_2360_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= AND_u32_u32_2360_inst_req_1;
      AND_u32_u32_2360_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAnd",
          name => "ApIntAnd_group_27",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00111111111111111111111110000000",
          constant_width => 32,
          buffering  => 1,
          flow_through => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 27
    -- shared split operator group (28) : AND_u32_u32_2508_inst 
    ApIntAnd_group_28: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= tmp10x_xix_xi30_2336;
      iNsTr_140_2509 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= AND_u32_u32_2508_inst_req_0;
      AND_u32_u32_2508_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= AND_u32_u32_2508_inst_req_1;
      AND_u32_u32_2508_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAnd",
          name => "ApIntAnd_group_28",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "10000000000000000000000000000000",
          constant_width => 32,
          buffering  => 1,
          flow_through => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 28
    -- shared split operator group (29) : AND_u32_u32_2514_inst 
    ApIntAnd_group_29: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= iNsTr_139_2503;
      iNsTr_141_2515 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= AND_u32_u32_2514_inst_req_0;
      AND_u32_u32_2514_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= AND_u32_u32_2514_inst_req_1;
      AND_u32_u32_2514_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAnd",
          name => "ApIntAnd_group_29",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000011111111",
          constant_width => 32,
          buffering  => 1,
          flow_through => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 29
    -- shared split operator group (30) : AND_u32_u32_2526_inst 
    ApIntAnd_group_30: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= xx_xlcssa19_2493;
      iNsTr_143_2527 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= AND_u32_u32_2526_inst_req_0;
      AND_u32_u32_2526_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= AND_u32_u32_2526_inst_req_1;
      AND_u32_u32_2526_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAnd",
          name => "ApIntAnd_group_30",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000100000000000000000000000",
          constant_width => 32,
          buffering  => 1,
          flow_through => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 30
    -- shared split operator group (31) : AND_u32_u32_2580_inst 
    ApIntAnd_group_31: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= iNsTr_206_2575;
      iNsTr_207_2581 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= AND_u32_u32_2580_inst_req_0;
      AND_u32_u32_2580_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= AND_u32_u32_2580_inst_req_1;
      AND_u32_u32_2580_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAnd",
          name => "ApIntAnd_group_31",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000100000000000000000000000",
          constant_width => 32,
          buffering  => 1,
          flow_through => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 31
    -- shared split operator group (32) : AND_u32_u32_2653_inst 
    ApIntAnd_group_32: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= tempx_x0x_xlcssax_xix_xi50_2642;
      iNsTr_177_2654 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= AND_u32_u32_2653_inst_req_0;
      AND_u32_u32_2653_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= AND_u32_u32_2653_inst_req_1;
      AND_u32_u32_2653_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAnd",
          name => "ApIntAnd_group_32",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000011111111111111111111111",
          constant_width => 32,
          buffering  => 1,
          flow_through => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 32
    -- shared split operator group (33) : AND_u32_u32_2734_inst 
    ApIntAnd_group_33: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= iNsTr_64_2729;
      iNsTr_65_2735 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= AND_u32_u32_2734_inst_req_0;
      AND_u32_u32_2734_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= AND_u32_u32_2734_inst_req_1;
      AND_u32_u32_2734_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAnd",
          name => "ApIntAnd_group_33",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000011111111",
          constant_width => 32,
          buffering  => 1,
          flow_through => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 33
    -- shared split operator group (34) : AND_u32_u32_2746_inst 
    ApIntAnd_group_34: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= iNsTr_66_2741;
      iNsTr_67_2747 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= AND_u32_u32_2746_inst_req_0;
      AND_u32_u32_2746_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= AND_u32_u32_2746_inst_req_1;
      AND_u32_u32_2746_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAnd",
          name => "ApIntAnd_group_34",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000011111111",
          constant_width => 32,
          buffering  => 1,
          flow_through => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 34
    -- shared split operator group (35) : AND_u32_u32_2758_inst 
    ApIntAnd_group_35: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= iNsTr_68_2753;
      iNsTr_69_2759 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= AND_u32_u32_2758_inst_req_0;
      AND_u32_u32_2758_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= AND_u32_u32_2758_inst_req_1;
      AND_u32_u32_2758_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAnd",
          name => "ApIntAnd_group_35",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00111111111111111111111110000000",
          constant_width => 32,
          buffering  => 1,
          flow_through => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 35
    -- shared split operator group (36) : AND_u32_u32_2776_inst 
    ApIntAnd_group_36: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= iNsTr_71_2771;
      iNsTr_72_2777 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= AND_u32_u32_2776_inst_req_0;
      AND_u32_u32_2776_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= AND_u32_u32_2776_inst_req_1;
      AND_u32_u32_2776_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAnd",
          name => "ApIntAnd_group_36",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000001111111111111111",
          constant_width => 32,
          buffering  => 1,
          flow_through => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 36
    -- shared split operator group (37) : AND_u32_u32_2793_inst 
    ApIntAnd_group_37: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= iNsTr_74_2788;
      iNsTr_75_2794 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= AND_u32_u32_2793_inst_req_0;
      AND_u32_u32_2793_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= AND_u32_u32_2793_inst_req_1;
      AND_u32_u32_2793_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAnd",
          name => "ApIntAnd_group_37",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "10000000000000000000000000000000",
          constant_width => 32,
          buffering  => 1,
          flow_through => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 37
    -- shared split operator group (38) : AND_u32_u32_2960_inst 
    ApIntAnd_group_38: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= tempx_x0x_xphx_xix_xi14_2949;
      iNsTr_104_2961 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= AND_u32_u32_2960_inst_req_0;
      AND_u32_u32_2960_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= AND_u32_u32_2960_inst_req_1;
      AND_u32_u32_2960_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAnd",
          name => "ApIntAnd_group_38",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000100000000000000000000000",
          constant_width => 32,
          buffering  => 1,
          flow_through => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 38
    -- shared split operator group (39) : AND_u32_u32_3014_inst 
    ApIntAnd_group_39: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= iNsTr_170_3009;
      iNsTr_171_3015 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= AND_u32_u32_3014_inst_req_0;
      AND_u32_u32_3014_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= AND_u32_u32_3014_inst_req_1;
      AND_u32_u32_3014_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAnd",
          name => "ApIntAnd_group_39",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000100000000000000000000000",
          constant_width => 32,
          buffering  => 1,
          flow_through => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 39
    -- shared split operator group (40) : AND_u32_u32_3092_inst 
    ApIntAnd_group_40: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= tempx_x0x_xlcssax_xix_xi26_3081;
      iNsTr_129_3093 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= AND_u32_u32_3092_inst_req_0;
      AND_u32_u32_3092_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= AND_u32_u32_3092_inst_req_1;
      AND_u32_u32_3092_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAnd",
          name => "ApIntAnd_group_40",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000011111111111111111111111",
          constant_width => 32,
          buffering  => 1,
          flow_through => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 40
    -- shared split operator group (41) : AND_u32_u32_3180_inst 
    ApIntAnd_group_41: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= iNsTr_88_3175;
      iNsTr_89_3181 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= AND_u32_u32_3180_inst_req_0;
      AND_u32_u32_3180_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= AND_u32_u32_3180_inst_req_1;
      AND_u32_u32_3180_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAnd",
          name => "ApIntAnd_group_41",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000011111111",
          constant_width => 32,
          buffering  => 1,
          flow_through => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 41
    -- shared split operator group (42) : AND_u32_u32_3192_inst 
    ApIntAnd_group_42: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= iNsTr_90_3187;
      iNsTr_91_3193 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= AND_u32_u32_3192_inst_req_0;
      AND_u32_u32_3192_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= AND_u32_u32_3192_inst_req_1;
      AND_u32_u32_3192_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAnd",
          name => "ApIntAnd_group_42",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000011111111",
          constant_width => 32,
          buffering  => 1,
          flow_through => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 42
    -- shared split operator group (43) : AND_u32_u32_3204_inst 
    ApIntAnd_group_43: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= iNsTr_92_3199;
      iNsTr_93_3205 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= AND_u32_u32_3204_inst_req_0;
      AND_u32_u32_3204_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= AND_u32_u32_3204_inst_req_1;
      AND_u32_u32_3204_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAnd",
          name => "ApIntAnd_group_43",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00111111111111111111111110000000",
          constant_width => 32,
          buffering  => 1,
          flow_through => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 43
    -- shared split operator group (44) : AND_u32_u32_3222_inst 
    ApIntAnd_group_44: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= iNsTr_95_3217;
      iNsTr_96_3223 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= AND_u32_u32_3222_inst_req_0;
      AND_u32_u32_3222_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= AND_u32_u32_3222_inst_req_1;
      AND_u32_u32_3222_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAnd",
          name => "ApIntAnd_group_44",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000001111111111111111",
          constant_width => 32,
          buffering  => 1,
          flow_through => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 44
    -- shared split operator group (45) : AND_u32_u32_3239_inst 
    ApIntAnd_group_45: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= iNsTr_98_3234;
      iNsTr_99_3240 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= AND_u32_u32_3239_inst_req_0;
      AND_u32_u32_3239_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= AND_u32_u32_3239_inst_req_1;
      AND_u32_u32_3239_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAnd",
          name => "ApIntAnd_group_45",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "10000000000000000000000000000000",
          constant_width => 32,
          buffering  => 1,
          flow_through => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 45
    -- shared split operator group (46) : AND_u32_u32_3406_inst 
    ApIntAnd_group_46: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= tempx_x0x_xphx_xix_xi_3395;
      iNsTr_121_3407 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= AND_u32_u32_3406_inst_req_0;
      AND_u32_u32_3406_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= AND_u32_u32_3406_inst_req_1;
      AND_u32_u32_3406_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAnd",
          name => "ApIntAnd_group_46",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000100000000000000000000000",
          constant_width => 32,
          buffering  => 1,
          flow_through => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 46
    -- shared split operator group (47) : AND_u32_u32_3460_inst 
    ApIntAnd_group_47: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= iNsTr_194_3455;
      iNsTr_195_3461 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= AND_u32_u32_3460_inst_req_0;
      AND_u32_u32_3460_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= AND_u32_u32_3460_inst_req_1;
      AND_u32_u32_3460_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAnd",
          name => "ApIntAnd_group_47",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000100000000000000000000000",
          constant_width => 32,
          buffering  => 1,
          flow_through => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 47
    -- shared split operator group (48) : AND_u32_u32_3538_inst 
    ApIntAnd_group_48: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= tempx_x0x_xlcssax_xix_xi_3527;
      iNsTr_158_3539 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= AND_u32_u32_3538_inst_req_0;
      AND_u32_u32_3538_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= AND_u32_u32_3538_inst_req_1;
      AND_u32_u32_3538_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAnd",
          name => "ApIntAnd_group_48",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000011111111111111111111111",
          constant_width => 32,
          buffering  => 1,
          flow_through => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 48
    -- shared split operator group (49) : AND_u32_u32_3712_inst 
    ApIntAnd_group_49: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= iNsTr_147_3707;
      iNsTr_148_3713 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= AND_u32_u32_3712_inst_req_0;
      AND_u32_u32_3712_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= AND_u32_u32_3712_inst_req_1;
      AND_u32_u32_3712_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAnd",
          name => "ApIntAnd_group_49",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00111111111111111111111110000000",
          constant_width => 32,
          buffering  => 1,
          flow_through => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 49
    -- shared split operator group (50) : AND_u32_u32_3860_inst 
    ApIntAnd_group_50: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= tmp10x_xi55_3701;
      iNsTr_239_3861 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= AND_u32_u32_3860_inst_req_0;
      AND_u32_u32_3860_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= AND_u32_u32_3860_inst_req_1;
      AND_u32_u32_3860_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAnd",
          name => "ApIntAnd_group_50",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "10000000000000000000000000000000",
          constant_width => 32,
          buffering  => 1,
          flow_through => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 50
    -- shared split operator group (51) : AND_u32_u32_3866_inst 
    ApIntAnd_group_51: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= iNsTr_238_3855;
      iNsTr_240_3867 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= AND_u32_u32_3866_inst_req_0;
      AND_u32_u32_3866_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= AND_u32_u32_3866_inst_req_1;
      AND_u32_u32_3866_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAnd",
          name => "ApIntAnd_group_51",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000011111111",
          constant_width => 32,
          buffering  => 1,
          flow_through => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 51
    -- shared split operator group (52) : AND_u32_u32_3878_inst 
    ApIntAnd_group_52: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= xx_xlcssa4_3845;
      iNsTr_242_3879 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= AND_u32_u32_3878_inst_req_0;
      AND_u32_u32_3878_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= AND_u32_u32_3878_inst_req_1;
      AND_u32_u32_3878_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAnd",
          name => "ApIntAnd_group_52",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000100000000000000000000000",
          constant_width => 32,
          buffering  => 1,
          flow_through => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 52
    -- shared split operator group (53) : AND_u32_u32_3932_inst 
    ApIntAnd_group_53: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= iNsTr_256_3927;
      iNsTr_257_3933 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= AND_u32_u32_3932_inst_req_0;
      AND_u32_u32_3932_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= AND_u32_u32_3932_inst_req_1;
      AND_u32_u32_3932_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAnd",
          name => "ApIntAnd_group_53",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000100000000000000000000000",
          constant_width => 32,
          buffering  => 1,
          flow_through => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 53
    -- shared split operator group (54) : AND_u32_u32_4005_inst 
    ApIntAnd_group_54: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= tempx_x0x_xlcssax_xi_3994;
      iNsTr_249_4006 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= AND_u32_u32_4005_inst_req_0;
      AND_u32_u32_4005_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= AND_u32_u32_4005_inst_req_1;
      AND_u32_u32_4005_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAnd",
          name => "ApIntAnd_group_54",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000011111111111111111111111",
          constant_width => 32,
          buffering  => 1,
          flow_through => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 54
    -- shared split operator group (55) : EQ_f32_u1_2341_inst 
    ApFloatUeq_group_55: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= iNsTr_32_2332;
      iNsTr_33_2342 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= EQ_f32_u1_2341_inst_req_0;
      EQ_f32_u1_2341_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= EQ_f32_u1_2341_inst_req_1;
      EQ_f32_u1_2341_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApFloatUeq",
          name => "ApFloatUeq_group_55",
          input1_is_int => false, 
          input1_characteristic_width => 8, 
          input1_mantissa_width    => 23, 
          iwidth_1  => 32,
          input2_is_int => false, 
          input2_characteristic_width => 8, 
          input2_mantissa_width => 23, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "00000000000000000000000000000000",
          constant_width => 32,
          buffering  => 1,
          flow_through => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 55
    -- shared split operator group (56) : EQ_f32_u1_2715_inst 
    ApFloatUeq_group_56: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= iNsTr_43_2696;
      iNsTr_45_2716 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= EQ_f32_u1_2715_inst_req_0;
      EQ_f32_u1_2715_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= EQ_f32_u1_2715_inst_req_1;
      EQ_f32_u1_2715_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApFloatUeq",
          name => "ApFloatUeq_group_56",
          input1_is_int => false, 
          input1_characteristic_width => 8, 
          input1_mantissa_width    => 23, 
          iwidth_1  => 32,
          input2_is_int => false, 
          input2_characteristic_width => 8, 
          input2_mantissa_width => 23, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "00000000000000000000000000000000",
          constant_width => 32,
          buffering  => 1,
          flow_through => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 56
    -- shared split operator group (57) : EQ_f32_u1_3161_inst 
    ApFloatUeq_group_57: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= torque_refx_x0_2190;
      iNsTr_62_3162 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= EQ_f32_u1_3161_inst_req_0;
      EQ_f32_u1_3161_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= EQ_f32_u1_3161_inst_req_1;
      EQ_f32_u1_3161_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApFloatUeq",
          name => "ApFloatUeq_group_57",
          input1_is_int => false, 
          input1_characteristic_width => 8, 
          input1_mantissa_width    => 23, 
          iwidth_1  => 32,
          input2_is_int => false, 
          input2_characteristic_width => 8, 
          input2_mantissa_width => 23, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "00000000000000000000000000000000",
          constant_width => 32,
          buffering  => 1,
          flow_through => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 57
    -- shared split operator group (58) : EQ_f32_u1_3678_inst 
    ApFloatUeq_group_58: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= iNsTr_114_3647;
      iNsTr_186_3679 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= EQ_f32_u1_3678_inst_req_0;
      EQ_f32_u1_3678_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= EQ_f32_u1_3678_inst_req_1;
      EQ_f32_u1_3678_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApFloatUeq",
          name => "ApFloatUeq_group_58",
          input1_is_int => false, 
          input1_characteristic_width => 8, 
          input1_mantissa_width    => 23, 
          iwidth_1  => 32,
          input2_is_int => false, 
          input2_characteristic_width => 8, 
          input2_mantissa_width => 23, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "00000000000000000000000000000000",
          constant_width => 32,
          buffering  => 1,
          flow_through => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 58
    -- shared split operator group (59) : EQ_u32_u1_2532_inst 
    ApIntEq_group_59: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= iNsTr_143_2527;
      iNsTr_144_2533 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= EQ_u32_u1_2532_inst_req_0;
      EQ_u32_u1_2532_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= EQ_u32_u1_2532_inst_req_1;
      EQ_u32_u1_2532_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntEq",
          name => "ApIntEq_group_59",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "00000000000000000000000000000000",
          constant_width => 32,
          buffering  => 1,
          flow_through => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 59
    -- shared split operator group (60) : EQ_u32_u1_2586_inst 
    ApIntEq_group_60: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= iNsTr_207_2581;
      iNsTr_208_2587 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= EQ_u32_u1_2586_inst_req_0;
      EQ_u32_u1_2586_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= EQ_u32_u1_2586_inst_req_1;
      EQ_u32_u1_2586_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntEq",
          name => "ApIntEq_group_60",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "00000000000000000000000000000000",
          constant_width => 32,
          buffering  => 1,
          flow_through => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 60
    -- shared split operator group (61) : EQ_u32_u1_2966_inst 
    ApIntEq_group_61: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= iNsTr_104_2961;
      iNsTr_105_2967 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= EQ_u32_u1_2966_inst_req_0;
      EQ_u32_u1_2966_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= EQ_u32_u1_2966_inst_req_1;
      EQ_u32_u1_2966_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntEq",
          name => "ApIntEq_group_61",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "00000000000000000000000000000000",
          constant_width => 32,
          buffering  => 1,
          flow_through => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 61
    -- shared split operator group (62) : EQ_u32_u1_3020_inst 
    ApIntEq_group_62: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= iNsTr_171_3015;
      iNsTr_172_3021 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= EQ_u32_u1_3020_inst_req_0;
      EQ_u32_u1_3020_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= EQ_u32_u1_3020_inst_req_1;
      EQ_u32_u1_3020_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntEq",
          name => "ApIntEq_group_62",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "00000000000000000000000000000000",
          constant_width => 32,
          buffering  => 1,
          flow_through => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 62
    -- shared split operator group (63) : EQ_u32_u1_3412_inst 
    ApIntEq_group_63: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= iNsTr_121_3407;
      iNsTr_122_3413 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= EQ_u32_u1_3412_inst_req_0;
      EQ_u32_u1_3412_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= EQ_u32_u1_3412_inst_req_1;
      EQ_u32_u1_3412_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntEq",
          name => "ApIntEq_group_63",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "00000000000000000000000000000000",
          constant_width => 32,
          buffering  => 1,
          flow_through => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 63
    -- shared split operator group (64) : EQ_u32_u1_3466_inst 
    ApIntEq_group_64: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= iNsTr_195_3461;
      iNsTr_196_3467 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= EQ_u32_u1_3466_inst_req_0;
      EQ_u32_u1_3466_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= EQ_u32_u1_3466_inst_req_1;
      EQ_u32_u1_3466_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntEq",
          name => "ApIntEq_group_64",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "00000000000000000000000000000000",
          constant_width => 32,
          buffering  => 1,
          flow_through => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 64
    -- shared split operator group (65) : EQ_u32_u1_3884_inst 
    ApIntEq_group_65: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= iNsTr_242_3879;
      iNsTr_243_3885 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= EQ_u32_u1_3884_inst_req_0;
      EQ_u32_u1_3884_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= EQ_u32_u1_3884_inst_req_1;
      EQ_u32_u1_3884_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntEq",
          name => "ApIntEq_group_65",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "00000000000000000000000000000000",
          constant_width => 32,
          buffering  => 1,
          flow_through => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 65
    -- shared split operator group (66) : EQ_u32_u1_3938_inst 
    ApIntEq_group_66: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= iNsTr_257_3933;
      iNsTr_258_3939 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= EQ_u32_u1_3938_inst_req_0;
      EQ_u32_u1_3938_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= EQ_u32_u1_3938_inst_req_1;
      EQ_u32_u1_3938_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntEq",
          name => "ApIntEq_group_66",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "00000000000000000000000000000000",
          constant_width => 32,
          buffering  => 1,
          flow_through => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 66
    -- shared split operator group (67) : LSHR_u32_u32_2388_inst 
    ApIntLSHR_group_67: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= xx_x016x_xix_xix_xi31_2370;
      iNsTr_78_2389 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= LSHR_u32_u32_2388_inst_req_0;
      LSHR_u32_u32_2388_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= LSHR_u32_u32_2388_inst_req_1;
      LSHR_u32_u32_2388_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntLSHR",
          name => "ApIntLSHR_group_67",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000001",
          constant_width => 32,
          buffering  => 1,
          flow_through => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 67
    -- shared split operator group (68) : LSHR_u32_u32_2502_inst 
    ApIntLSHR_group_68: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= tmp10x_xix_xi30_2336;
      iNsTr_139_2503 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= LSHR_u32_u32_2502_inst_req_0;
      LSHR_u32_u32_2502_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= LSHR_u32_u32_2502_inst_req_1;
      LSHR_u32_u32_2502_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntLSHR",
          name => "ApIntLSHR_group_68",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000010111",
          constant_width => 32,
          buffering  => 1,
          flow_through => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 68
    -- shared split operator group (69) : LSHR_u32_u32_2728_inst 
    ApIntLSHR_group_69: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= tmp10x_xix_xi1_2706;
      iNsTr_64_2729 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= LSHR_u32_u32_2728_inst_req_0;
      LSHR_u32_u32_2728_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= LSHR_u32_u32_2728_inst_req_1;
      LSHR_u32_u32_2728_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntLSHR",
          name => "ApIntLSHR_group_69",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000010111",
          constant_width => 32,
          buffering  => 1,
          flow_through => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 69
    -- shared split operator group (70) : LSHR_u32_u32_2740_inst 
    ApIntLSHR_group_70: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= tmp6x_xix_xi2_2710;
      iNsTr_66_2741 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= LSHR_u32_u32_2740_inst_req_0;
      LSHR_u32_u32_2740_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= LSHR_u32_u32_2740_inst_req_1;
      LSHR_u32_u32_2740_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntLSHR",
          name => "ApIntLSHR_group_70",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000010111",
          constant_width => 32,
          buffering  => 1,
          flow_through => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 70
    -- shared split operator group (71) : LSHR_u32_u32_2770_inst 
    ApIntLSHR_group_71: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= tmp6x_xix_xi2_2710;
      iNsTr_71_2771 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= LSHR_u32_u32_2770_inst_req_0;
      LSHR_u32_u32_2770_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= LSHR_u32_u32_2770_inst_req_1;
      LSHR_u32_u32_2770_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntLSHR",
          name => "ApIntLSHR_group_71",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000111",
          constant_width => 32,
          buffering  => 1,
          flow_through => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 71
    -- shared split operator group (72) : LSHR_u32_u32_2831_inst 
    ApIntLSHR_group_72: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= xx_x016x_xix_xix_xi3_2813;
      iNsTr_125_2832 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= LSHR_u32_u32_2831_inst_req_0;
      LSHR_u32_u32_2831_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= LSHR_u32_u32_2831_inst_req_1;
      LSHR_u32_u32_2831_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntLSHR",
          name => "ApIntLSHR_group_72",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000001",
          constant_width => 32,
          buffering  => 1,
          flow_through => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 72
    -- shared split operator group (73) : LSHR_u32_u32_3174_inst 
    ApIntLSHR_group_73: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= tmp10x_xix_xi_3145;
      iNsTr_88_3175 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= LSHR_u32_u32_3174_inst_req_0;
      LSHR_u32_u32_3174_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= LSHR_u32_u32_3174_inst_req_1;
      LSHR_u32_u32_3174_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntLSHR",
          name => "ApIntLSHR_group_73",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000010111",
          constant_width => 32,
          buffering  => 1,
          flow_through => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 73
    -- shared split operator group (74) : LSHR_u32_u32_3186_inst 
    ApIntLSHR_group_74: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= tmp6x_xix_xi_3156;
      iNsTr_90_3187 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= LSHR_u32_u32_3186_inst_req_0;
      LSHR_u32_u32_3186_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= LSHR_u32_u32_3186_inst_req_1;
      LSHR_u32_u32_3186_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntLSHR",
          name => "ApIntLSHR_group_74",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000010111",
          constant_width => 32,
          buffering  => 1,
          flow_through => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 74
    -- shared split operator group (75) : LSHR_u32_u32_3216_inst 
    ApIntLSHR_group_75: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= tmp6x_xix_xi_3156;
      iNsTr_95_3217 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= LSHR_u32_u32_3216_inst_req_0;
      LSHR_u32_u32_3216_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= LSHR_u32_u32_3216_inst_req_1;
      LSHR_u32_u32_3216_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntLSHR",
          name => "ApIntLSHR_group_75",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000111",
          constant_width => 32,
          buffering  => 1,
          flow_through => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 75
    -- shared split operator group (76) : LSHR_u32_u32_3277_inst 
    ApIntLSHR_group_76: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= xx_x016x_xix_xix_xi_3259;
      iNsTr_154_3278 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= LSHR_u32_u32_3277_inst_req_0;
      LSHR_u32_u32_3277_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= LSHR_u32_u32_3277_inst_req_1;
      LSHR_u32_u32_3277_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntLSHR",
          name => "ApIntLSHR_group_76",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000001",
          constant_width => 32,
          buffering  => 1,
          flow_through => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 76
    -- shared split operator group (77) : LSHR_u32_u32_3740_inst 
    ApIntLSHR_group_77: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= xx_x016x_xix_xi_3722;
      iNsTr_183_3741 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= LSHR_u32_u32_3740_inst_req_0;
      LSHR_u32_u32_3740_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= LSHR_u32_u32_3740_inst_req_1;
      LSHR_u32_u32_3740_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntLSHR",
          name => "ApIntLSHR_group_77",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000001",
          constant_width => 32,
          buffering  => 1,
          flow_through => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 77
    -- shared split operator group (78) : LSHR_u32_u32_3854_inst 
    ApIntLSHR_group_78: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= tmp10x_xi55_3701;
      iNsTr_238_3855 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= LSHR_u32_u32_3854_inst_req_0;
      LSHR_u32_u32_3854_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= LSHR_u32_u32_3854_inst_req_1;
      LSHR_u32_u32_3854_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntLSHR",
          name => "ApIntLSHR_group_78",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000010111",
          constant_width => 32,
          buffering  => 1,
          flow_through => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 78
    -- shared split operator group (79) : MUL_f32_f32_2320_inst MUL_f32_f32_2247_inst MUL_f32_f32_2099_inst MUL_f32_f32_2088_inst MUL_f32_f32_2149_inst MUL_f32_f32_2186_inst MUL_f32_f32_2235_inst MUL_f32_f32_2268_inst MUL_f32_f32_2300_inst MUL_f32_f32_2280_inst MUL_f32_f32_2326_inst MUL_f32_f32_2288_inst MUL_f32_f32_2695_inst MUL_f32_f32_2701_inst MUL_f32_f32_3140_inst MUL_f32_f32_3585_inst MUL_f32_f32_3596_inst MUL_f32_f32_3641_inst 
    ApFloatMul_group_79: Block -- 
      signal data_in: std_logic_vector(1151 downto 0);
      signal data_out: std_logic_vector(575 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 17 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 17 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 17 downto 0);
      signal guard_vector : std_logic_vector( 17 downto 0);
      constant inBUFs : IntegerArray(17 downto 0) := (17 => 1, 16 => 1, 15 => 1, 14 => 1, 13 => 1, 12 => 1, 11 => 1, 10 => 1, 9 => 1, 8 => 1, 7 => 1, 6 => 1, 5 => 1, 4 => 1, 3 => 1, 2 => 1, 1 => 1, 0 => 1);
      constant outBUFs : IntegerArray(17 downto 0) := (17 => 1, 16 => 1, 15 => 1, 14 => 1, 13 => 1, 12 => 1, 11 => 1, 10 => 1, 9 => 1, 8 => 1, 7 => 1, 6 => 1, 5 => 1, 4 => 1, 3 => 1, 2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(17 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false, 8 => false, 9 => false, 10 => false, 11 => false, 12 => false, 13 => false, 14 => false, 15 => false, 16 => false, 17 => false);
      constant guardBuffering: IntegerArray(17 downto 0)  := (0 => 1, 1 => 1, 2 => 1, 3 => 1, 4 => 1, 5 => 1, 6 => 1, 7 => 1, 8 => 1, 9 => 1, 10 => 1, 11 => 1, 12 => 1, 13 => 1, 14 => 1, 15 => 1, 16 => 1, 17 => 1);
      -- 
    begin -- 
      data_in <= iNsTr_2_2069 & type_cast_2319_wire_constant & iNsTr_39_2242 & type_cast_2246_wire_constant & iNsTr_11_2094 & type_cast_2098_wire_constant & iNsTr_9_2083 & type_cast_2087_wire_constant & iNsTr_9_2083 & type_cast_2148_wire_constant & iNsTr_17_2155 & type_cast_2185_wire_constant & iNsTr_8_2078 & type_cast_2234_wire_constant & iNsTr_8_2078 & type_cast_2267_wire_constant & iNsTr_52_2295 & type_cast_2299_wire_constant & iNsTr_56_2275 & type_cast_2279_wire_constant & flux_rotor_prevx_x0_2045 & type_cast_2325_wire_constant & iNsTr_8_2078 & type_cast_2287_wire_constant & iNsTr_4_2072 & type_cast_2694_wire_constant & iNsTr_42_2683 & type_cast_2700_wire_constant & iNsTr_42_2683 & type_cast_3139_wire_constant & iNsTr_82_3580 & type_cast_3584_wire_constant & iNsTr_84_3591 & type_cast_3595_wire_constant & iNsTr_82_3580 & type_cast_3640_wire_constant;
      iNsTr_30_2321 <= data_out(575 downto 544);
      iNsTr_40_2248 <= data_out(543 downto 512);
      iNsTr_12_2100 <= data_out(511 downto 480);
      iNsTr_10_2089 <= data_out(479 downto 448);
      iNsTr_16_2150 <= data_out(447 downto 416);
      phitmp_2187 <= data_out(415 downto 384);
      iNsTr_38_2236 <= data_out(383 downto 352);
      iNsTr_55_2269 <= data_out(351 downto 320);
      iNsTr_53_2301 <= data_out(319 downto 288);
      iNsTr_57_2281 <= data_out(287 downto 256);
      iNsTr_31_2327 <= data_out(255 downto 224);
      iNsTr_51_2289 <= data_out(223 downto 192);
      iNsTr_43_2696 <= data_out(191 downto 160);
      iNsTr_44_2702 <= data_out(159 downto 128);
      xx_xop_3141 <= data_out(127 downto 96);
      iNsTr_83_3586 <= data_out(95 downto 64);
      iNsTr_85_3597 <= data_out(63 downto 32);
      iNsTr_113_3642 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      guard_vector(8)  <=  '1';
      guard_vector(9)  <=  '1';
      guard_vector(10)  <=  '1';
      guard_vector(11)  <=  '1';
      guard_vector(12)  <=  '1';
      guard_vector(13)  <=  '1';
      guard_vector(14)  <=  '1';
      guard_vector(15)  <=  '1';
      guard_vector(16)  <=  '1';
      guard_vector(17)  <=  '1';
      reqL_unguarded(17) <= MUL_f32_f32_2320_inst_req_0;
      reqL_unguarded(16) <= MUL_f32_f32_2247_inst_req_0;
      reqL_unguarded(15) <= MUL_f32_f32_2099_inst_req_0;
      reqL_unguarded(14) <= MUL_f32_f32_2088_inst_req_0;
      reqL_unguarded(13) <= MUL_f32_f32_2149_inst_req_0;
      reqL_unguarded(12) <= MUL_f32_f32_2186_inst_req_0;
      reqL_unguarded(11) <= MUL_f32_f32_2235_inst_req_0;
      reqL_unguarded(10) <= MUL_f32_f32_2268_inst_req_0;
      reqL_unguarded(9) <= MUL_f32_f32_2300_inst_req_0;
      reqL_unguarded(8) <= MUL_f32_f32_2280_inst_req_0;
      reqL_unguarded(7) <= MUL_f32_f32_2326_inst_req_0;
      reqL_unguarded(6) <= MUL_f32_f32_2288_inst_req_0;
      reqL_unguarded(5) <= MUL_f32_f32_2695_inst_req_0;
      reqL_unguarded(4) <= MUL_f32_f32_2701_inst_req_0;
      reqL_unguarded(3) <= MUL_f32_f32_3140_inst_req_0;
      reqL_unguarded(2) <= MUL_f32_f32_3585_inst_req_0;
      reqL_unguarded(1) <= MUL_f32_f32_3596_inst_req_0;
      reqL_unguarded(0) <= MUL_f32_f32_3641_inst_req_0;
      MUL_f32_f32_2320_inst_ack_0 <= ackL_unguarded(17);
      MUL_f32_f32_2247_inst_ack_0 <= ackL_unguarded(16);
      MUL_f32_f32_2099_inst_ack_0 <= ackL_unguarded(15);
      MUL_f32_f32_2088_inst_ack_0 <= ackL_unguarded(14);
      MUL_f32_f32_2149_inst_ack_0 <= ackL_unguarded(13);
      MUL_f32_f32_2186_inst_ack_0 <= ackL_unguarded(12);
      MUL_f32_f32_2235_inst_ack_0 <= ackL_unguarded(11);
      MUL_f32_f32_2268_inst_ack_0 <= ackL_unguarded(10);
      MUL_f32_f32_2300_inst_ack_0 <= ackL_unguarded(9);
      MUL_f32_f32_2280_inst_ack_0 <= ackL_unguarded(8);
      MUL_f32_f32_2326_inst_ack_0 <= ackL_unguarded(7);
      MUL_f32_f32_2288_inst_ack_0 <= ackL_unguarded(6);
      MUL_f32_f32_2695_inst_ack_0 <= ackL_unguarded(5);
      MUL_f32_f32_2701_inst_ack_0 <= ackL_unguarded(4);
      MUL_f32_f32_3140_inst_ack_0 <= ackL_unguarded(3);
      MUL_f32_f32_3585_inst_ack_0 <= ackL_unguarded(2);
      MUL_f32_f32_3596_inst_ack_0 <= ackL_unguarded(1);
      MUL_f32_f32_3641_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(17) <= MUL_f32_f32_2320_inst_req_1;
      reqR_unguarded(16) <= MUL_f32_f32_2247_inst_req_1;
      reqR_unguarded(15) <= MUL_f32_f32_2099_inst_req_1;
      reqR_unguarded(14) <= MUL_f32_f32_2088_inst_req_1;
      reqR_unguarded(13) <= MUL_f32_f32_2149_inst_req_1;
      reqR_unguarded(12) <= MUL_f32_f32_2186_inst_req_1;
      reqR_unguarded(11) <= MUL_f32_f32_2235_inst_req_1;
      reqR_unguarded(10) <= MUL_f32_f32_2268_inst_req_1;
      reqR_unguarded(9) <= MUL_f32_f32_2300_inst_req_1;
      reqR_unguarded(8) <= MUL_f32_f32_2280_inst_req_1;
      reqR_unguarded(7) <= MUL_f32_f32_2326_inst_req_1;
      reqR_unguarded(6) <= MUL_f32_f32_2288_inst_req_1;
      reqR_unguarded(5) <= MUL_f32_f32_2695_inst_req_1;
      reqR_unguarded(4) <= MUL_f32_f32_2701_inst_req_1;
      reqR_unguarded(3) <= MUL_f32_f32_3140_inst_req_1;
      reqR_unguarded(2) <= MUL_f32_f32_3585_inst_req_1;
      reqR_unguarded(1) <= MUL_f32_f32_3596_inst_req_1;
      reqR_unguarded(0) <= MUL_f32_f32_3641_inst_req_1;
      MUL_f32_f32_2320_inst_ack_1 <= ackR_unguarded(17);
      MUL_f32_f32_2247_inst_ack_1 <= ackR_unguarded(16);
      MUL_f32_f32_2099_inst_ack_1 <= ackR_unguarded(15);
      MUL_f32_f32_2088_inst_ack_1 <= ackR_unguarded(14);
      MUL_f32_f32_2149_inst_ack_1 <= ackR_unguarded(13);
      MUL_f32_f32_2186_inst_ack_1 <= ackR_unguarded(12);
      MUL_f32_f32_2235_inst_ack_1 <= ackR_unguarded(11);
      MUL_f32_f32_2268_inst_ack_1 <= ackR_unguarded(10);
      MUL_f32_f32_2300_inst_ack_1 <= ackR_unguarded(9);
      MUL_f32_f32_2280_inst_ack_1 <= ackR_unguarded(8);
      MUL_f32_f32_2326_inst_ack_1 <= ackR_unguarded(7);
      MUL_f32_f32_2288_inst_ack_1 <= ackR_unguarded(6);
      MUL_f32_f32_2695_inst_ack_1 <= ackR_unguarded(5);
      MUL_f32_f32_2701_inst_ack_1 <= ackR_unguarded(4);
      MUL_f32_f32_3140_inst_ack_1 <= ackR_unguarded(3);
      MUL_f32_f32_3585_inst_ack_1 <= ackR_unguarded(2);
      MUL_f32_f32_3596_inst_ack_1 <= ackR_unguarded(1);
      MUL_f32_f32_3641_inst_ack_1 <= ackR_unguarded(0);
      ApFloatMul_group_79_accessRegulator_0: access_regulator_base generic map (name => "ApFloatMul_group_79_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      ApFloatMul_group_79_accessRegulator_1: access_regulator_base generic map (name => "ApFloatMul_group_79_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      ApFloatMul_group_79_accessRegulator_2: access_regulator_base generic map (name => "ApFloatMul_group_79_accessRegulator_2", num_slots => 1) -- 
        port map (req => reqL_unregulated(2), -- 
          ack => ackL_unregulated(2),
          regulated_req => reqL(2),
          regulated_ack => ackL(2),
          release_req => reqR(2),
          release_ack => ackR(2),
          clk => clk, reset => reset); -- 
      ApFloatMul_group_79_accessRegulator_3: access_regulator_base generic map (name => "ApFloatMul_group_79_accessRegulator_3", num_slots => 1) -- 
        port map (req => reqL_unregulated(3), -- 
          ack => ackL_unregulated(3),
          regulated_req => reqL(3),
          regulated_ack => ackL(3),
          release_req => reqR(3),
          release_ack => ackR(3),
          clk => clk, reset => reset); -- 
      ApFloatMul_group_79_accessRegulator_4: access_regulator_base generic map (name => "ApFloatMul_group_79_accessRegulator_4", num_slots => 1) -- 
        port map (req => reqL_unregulated(4), -- 
          ack => ackL_unregulated(4),
          regulated_req => reqL(4),
          regulated_ack => ackL(4),
          release_req => reqR(4),
          release_ack => ackR(4),
          clk => clk, reset => reset); -- 
      ApFloatMul_group_79_accessRegulator_5: access_regulator_base generic map (name => "ApFloatMul_group_79_accessRegulator_5", num_slots => 1) -- 
        port map (req => reqL_unregulated(5), -- 
          ack => ackL_unregulated(5),
          regulated_req => reqL(5),
          regulated_ack => ackL(5),
          release_req => reqR(5),
          release_ack => ackR(5),
          clk => clk, reset => reset); -- 
      ApFloatMul_group_79_accessRegulator_6: access_regulator_base generic map (name => "ApFloatMul_group_79_accessRegulator_6", num_slots => 1) -- 
        port map (req => reqL_unregulated(6), -- 
          ack => ackL_unregulated(6),
          regulated_req => reqL(6),
          regulated_ack => ackL(6),
          release_req => reqR(6),
          release_ack => ackR(6),
          clk => clk, reset => reset); -- 
      ApFloatMul_group_79_accessRegulator_7: access_regulator_base generic map (name => "ApFloatMul_group_79_accessRegulator_7", num_slots => 1) -- 
        port map (req => reqL_unregulated(7), -- 
          ack => ackL_unregulated(7),
          regulated_req => reqL(7),
          regulated_ack => ackL(7),
          release_req => reqR(7),
          release_ack => ackR(7),
          clk => clk, reset => reset); -- 
      ApFloatMul_group_79_accessRegulator_8: access_regulator_base generic map (name => "ApFloatMul_group_79_accessRegulator_8", num_slots => 1) -- 
        port map (req => reqL_unregulated(8), -- 
          ack => ackL_unregulated(8),
          regulated_req => reqL(8),
          regulated_ack => ackL(8),
          release_req => reqR(8),
          release_ack => ackR(8),
          clk => clk, reset => reset); -- 
      ApFloatMul_group_79_accessRegulator_9: access_regulator_base generic map (name => "ApFloatMul_group_79_accessRegulator_9", num_slots => 1) -- 
        port map (req => reqL_unregulated(9), -- 
          ack => ackL_unregulated(9),
          regulated_req => reqL(9),
          regulated_ack => ackL(9),
          release_req => reqR(9),
          release_ack => ackR(9),
          clk => clk, reset => reset); -- 
      ApFloatMul_group_79_accessRegulator_10: access_regulator_base generic map (name => "ApFloatMul_group_79_accessRegulator_10", num_slots => 1) -- 
        port map (req => reqL_unregulated(10), -- 
          ack => ackL_unregulated(10),
          regulated_req => reqL(10),
          regulated_ack => ackL(10),
          release_req => reqR(10),
          release_ack => ackR(10),
          clk => clk, reset => reset); -- 
      ApFloatMul_group_79_accessRegulator_11: access_regulator_base generic map (name => "ApFloatMul_group_79_accessRegulator_11", num_slots => 1) -- 
        port map (req => reqL_unregulated(11), -- 
          ack => ackL_unregulated(11),
          regulated_req => reqL(11),
          regulated_ack => ackL(11),
          release_req => reqR(11),
          release_ack => ackR(11),
          clk => clk, reset => reset); -- 
      ApFloatMul_group_79_accessRegulator_12: access_regulator_base generic map (name => "ApFloatMul_group_79_accessRegulator_12", num_slots => 1) -- 
        port map (req => reqL_unregulated(12), -- 
          ack => ackL_unregulated(12),
          regulated_req => reqL(12),
          regulated_ack => ackL(12),
          release_req => reqR(12),
          release_ack => ackR(12),
          clk => clk, reset => reset); -- 
      ApFloatMul_group_79_accessRegulator_13: access_regulator_base generic map (name => "ApFloatMul_group_79_accessRegulator_13", num_slots => 1) -- 
        port map (req => reqL_unregulated(13), -- 
          ack => ackL_unregulated(13),
          regulated_req => reqL(13),
          regulated_ack => ackL(13),
          release_req => reqR(13),
          release_ack => ackR(13),
          clk => clk, reset => reset); -- 
      ApFloatMul_group_79_accessRegulator_14: access_regulator_base generic map (name => "ApFloatMul_group_79_accessRegulator_14", num_slots => 1) -- 
        port map (req => reqL_unregulated(14), -- 
          ack => ackL_unregulated(14),
          regulated_req => reqL(14),
          regulated_ack => ackL(14),
          release_req => reqR(14),
          release_ack => ackR(14),
          clk => clk, reset => reset); -- 
      ApFloatMul_group_79_accessRegulator_15: access_regulator_base generic map (name => "ApFloatMul_group_79_accessRegulator_15", num_slots => 1) -- 
        port map (req => reqL_unregulated(15), -- 
          ack => ackL_unregulated(15),
          regulated_req => reqL(15),
          regulated_ack => ackL(15),
          release_req => reqR(15),
          release_ack => ackR(15),
          clk => clk, reset => reset); -- 
      ApFloatMul_group_79_accessRegulator_16: access_regulator_base generic map (name => "ApFloatMul_group_79_accessRegulator_16", num_slots => 1) -- 
        port map (req => reqL_unregulated(16), -- 
          ack => ackL_unregulated(16),
          regulated_req => reqL(16),
          regulated_ack => ackL(16),
          release_req => reqR(16),
          release_ack => ackR(16),
          clk => clk, reset => reset); -- 
      ApFloatMul_group_79_accessRegulator_17: access_regulator_base generic map (name => "ApFloatMul_group_79_accessRegulator_17", num_slots => 1) -- 
        port map (req => reqL_unregulated(17), -- 
          ack => ackL_unregulated(17),
          regulated_req => reqL(17),
          regulated_ack => ackL(17),
          release_req => reqR(17),
          release_ack => ackR(17),
          clk => clk, reset => reset); -- 
      gI: SplitGuardInterface generic map(nreqs => 18, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      PipedFpOp: PipelinedFPOperator -- 
        generic map( -- 
          name => "ApFloatMul_group_79",
          operator_id => "ApFloatMul",
          exponent_width => 8,
          fraction_width => 23, 
          no_arbitration => false,
          num_reqs => 18,
          use_input_buffering => true,
          detailed_buffering_per_input => inBUFs,
          detailed_buffering_per_output => outBUFs -- 
        )
        port map ( reqL => reqL , ackL => ackL, reqR => reqR, ackR => ackR, dataL => data_in, dataR => data_out, clk => clk, reset => reset); -- 
      -- 
    end Block; -- split operator group 79
    -- shared split operator group (80) : NEQ_i32_u1_2540_inst 
    ApIntNe_group_80: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= type_cast_2536_wire;
      iNsTr_145_2541 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= NEQ_i32_u1_2540_inst_req_0;
      NEQ_i32_u1_2540_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= NEQ_i32_u1_2540_inst_req_1;
      NEQ_i32_u1_2540_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntNe",
          name => "ApIntNe_group_80",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "00000000000000000000000000000000",
          constant_width => 32,
          buffering  => 1,
          flow_through => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 80
    -- shared split operator group (81) : NEQ_i32_u1_2594_inst 
    ApIntNe_group_81: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= type_cast_2590_wire;
      iNsTr_209_2595 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= NEQ_i32_u1_2594_inst_req_0;
      NEQ_i32_u1_2594_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= NEQ_i32_u1_2594_inst_req_1;
      NEQ_i32_u1_2594_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntNe",
          name => "ApIntNe_group_81",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "00000000000000000000000000000000",
          constant_width => 32,
          buffering  => 1,
          flow_through => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 81
    -- shared split operator group (82) : NEQ_i32_u1_2974_inst 
    ApIntNe_group_82: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= type_cast_2970_wire;
      iNsTr_106_2975 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= NEQ_i32_u1_2974_inst_req_0;
      NEQ_i32_u1_2974_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= NEQ_i32_u1_2974_inst_req_1;
      NEQ_i32_u1_2974_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntNe",
          name => "ApIntNe_group_82",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "00000000000000000000000000000000",
          constant_width => 32,
          buffering  => 1,
          flow_through => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 82
    -- shared split operator group (83) : NEQ_i32_u1_3028_inst 
    ApIntNe_group_83: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= type_cast_3024_wire;
      iNsTr_173_3029 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= NEQ_i32_u1_3028_inst_req_0;
      NEQ_i32_u1_3028_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= NEQ_i32_u1_3028_inst_req_1;
      NEQ_i32_u1_3028_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntNe",
          name => "ApIntNe_group_83",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "00000000000000000000000000000000",
          constant_width => 32,
          buffering  => 1,
          flow_through => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 83
    -- shared split operator group (84) : NEQ_i32_u1_3420_inst 
    ApIntNe_group_84: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= type_cast_3416_wire;
      iNsTr_123_3421 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= NEQ_i32_u1_3420_inst_req_0;
      NEQ_i32_u1_3420_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= NEQ_i32_u1_3420_inst_req_1;
      NEQ_i32_u1_3420_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntNe",
          name => "ApIntNe_group_84",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "00000000000000000000000000000000",
          constant_width => 32,
          buffering  => 1,
          flow_through => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 84
    -- shared split operator group (85) : NEQ_i32_u1_3474_inst 
    ApIntNe_group_85: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= type_cast_3470_wire;
      iNsTr_197_3475 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= NEQ_i32_u1_3474_inst_req_0;
      NEQ_i32_u1_3474_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= NEQ_i32_u1_3474_inst_req_1;
      NEQ_i32_u1_3474_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntNe",
          name => "ApIntNe_group_85",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "00000000000000000000000000000000",
          constant_width => 32,
          buffering  => 1,
          flow_through => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 85
    -- shared split operator group (86) : NEQ_i32_u1_3892_inst 
    ApIntNe_group_86: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= type_cast_3888_wire;
      iNsTr_244_3893 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= NEQ_i32_u1_3892_inst_req_0;
      NEQ_i32_u1_3892_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= NEQ_i32_u1_3892_inst_req_1;
      NEQ_i32_u1_3892_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntNe",
          name => "ApIntNe_group_86",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "00000000000000000000000000000000",
          constant_width => 32,
          buffering  => 1,
          flow_through => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 86
    -- shared split operator group (87) : NEQ_i32_u1_3946_inst 
    ApIntNe_group_87: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= type_cast_3942_wire;
      iNsTr_259_3947 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= NEQ_i32_u1_3946_inst_req_0;
      NEQ_i32_u1_3946_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= NEQ_i32_u1_3946_inst_req_1;
      NEQ_i32_u1_3946_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntNe",
          name => "ApIntNe_group_87",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "00000000000000000000000000000000",
          constant_width => 32,
          buffering  => 1,
          flow_through => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 87
    -- shared split operator group (88) : OR_u32_u32_2366_inst 
    ApIntOr_group_88: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= iNsTr_48_2361;
      iNsTr_49_2367 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= OR_u32_u32_2366_inst_req_0;
      OR_u32_u32_2366_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= OR_u32_u32_2366_inst_req_1;
      OR_u32_u32_2366_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntOr",
          name => "ApIntOr_group_88",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "01000000000000000000000000000000",
          constant_width => 32,
          buffering  => 1,
          flow_through => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 88
    -- shared split operator group (89) : OR_u32_u32_2670_inst 
    ApIntOr_group_89: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= iNsTr_177_2654 & iNsTr_140_2509;
      iNsTr_180_2671 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= OR_u32_u32_2670_inst_req_0;
      OR_u32_u32_2670_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= OR_u32_u32_2670_inst_req_1;
      OR_u32_u32_2670_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntOr",
          name => "ApIntOr_group_89",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 89
    -- shared split operator group (90) : OR_u32_u32_2675_inst 
    ApIntOr_group_90: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= iNsTr_180_2671 & iNsTr_179_2666;
      iNsTr_181_2676 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= OR_u32_u32_2675_inst_req_0;
      OR_u32_u32_2675_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= OR_u32_u32_2675_inst_req_1;
      OR_u32_u32_2675_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntOr",
          name => "ApIntOr_group_90",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 90
    -- shared split operator group (91) : OR_u32_u32_2764_inst 
    ApIntOr_group_91: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= iNsTr_69_2759;
      iNsTr_70_2765 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= OR_u32_u32_2764_inst_req_0;
      OR_u32_u32_2764_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= OR_u32_u32_2764_inst_req_1;
      OR_u32_u32_2764_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntOr",
          name => "ApIntOr_group_91",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "01000000000000000000000000000000",
          constant_width => 32,
          buffering  => 1,
          flow_through => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 91
    -- shared split operator group (92) : OR_u32_u32_2782_inst 
    ApIntOr_group_92: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= iNsTr_72_2777;
      iNsTr_73_2783 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= OR_u32_u32_2782_inst_req_0;
      OR_u32_u32_2782_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= OR_u32_u32_2782_inst_req_1;
      OR_u32_u32_2782_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntOr",
          name => "ApIntOr_group_92",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000010000000000000000",
          constant_width => 32,
          buffering  => 1,
          flow_through => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 92
    -- shared split operator group (93) : OR_u32_u32_3109_inst 
    ApIntOr_group_93: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= iNsTr_129_3093 & iNsTr_75_2794;
      iNsTr_132_3110 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= OR_u32_u32_3109_inst_req_0;
      OR_u32_u32_3109_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= OR_u32_u32_3109_inst_req_1;
      OR_u32_u32_3109_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntOr",
          name => "ApIntOr_group_93",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 93
    -- shared split operator group (94) : OR_u32_u32_3114_inst 
    ApIntOr_group_94: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= iNsTr_132_3110 & iNsTr_131_3105;
      iNsTr_133_3115 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= OR_u32_u32_3114_inst_req_0;
      OR_u32_u32_3114_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= OR_u32_u32_3114_inst_req_1;
      OR_u32_u32_3114_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntOr",
          name => "ApIntOr_group_94",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 94
    -- shared split operator group (95) : OR_u32_u32_3210_inst 
    ApIntOr_group_95: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= iNsTr_93_3205;
      iNsTr_94_3211 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= OR_u32_u32_3210_inst_req_0;
      OR_u32_u32_3210_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= OR_u32_u32_3210_inst_req_1;
      OR_u32_u32_3210_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntOr",
          name => "ApIntOr_group_95",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "01000000000000000000000000000000",
          constant_width => 32,
          buffering  => 1,
          flow_through => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 95
    -- shared split operator group (96) : OR_u32_u32_3228_inst 
    ApIntOr_group_96: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= iNsTr_96_3223;
      iNsTr_97_3229 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= OR_u32_u32_3228_inst_req_0;
      OR_u32_u32_3228_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= OR_u32_u32_3228_inst_req_1;
      OR_u32_u32_3228_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntOr",
          name => "ApIntOr_group_96",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000010000000000000000",
          constant_width => 32,
          buffering  => 1,
          flow_through => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 96
    -- shared split operator group (97) : OR_u32_u32_3555_inst 
    ApIntOr_group_97: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= iNsTr_158_3539 & iNsTr_99_3240;
      iNsTr_161_3556 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= OR_u32_u32_3555_inst_req_0;
      OR_u32_u32_3555_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= OR_u32_u32_3555_inst_req_1;
      OR_u32_u32_3555_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntOr",
          name => "ApIntOr_group_97",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 97
    -- shared split operator group (98) : OR_u32_u32_3560_inst 
    ApIntOr_group_98: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= iNsTr_161_3556 & iNsTr_160_3551;
      iNsTr_162_3561 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= OR_u32_u32_3560_inst_req_0;
      OR_u32_u32_3560_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= OR_u32_u32_3560_inst_req_1;
      OR_u32_u32_3560_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntOr",
          name => "ApIntOr_group_98",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 98
    -- shared split operator group (99) : OR_u32_u32_3718_inst 
    ApIntOr_group_99: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= iNsTr_148_3713;
      iNsTr_149_3719 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= OR_u32_u32_3718_inst_req_0;
      OR_u32_u32_3718_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= OR_u32_u32_3718_inst_req_1;
      OR_u32_u32_3718_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntOr",
          name => "ApIntOr_group_99",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "01000000000000000000000000000000",
          constant_width => 32,
          buffering  => 1,
          flow_through => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 99
    -- shared split operator group (100) : OR_u32_u32_4022_inst 
    ApIntOr_group_100: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= iNsTr_251_4018 & iNsTr_239_3861;
      iNsTr_252_4023 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= OR_u32_u32_4022_inst_req_0;
      OR_u32_u32_4022_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= OR_u32_u32_4022_inst_req_1;
      OR_u32_u32_4022_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntOr",
          name => "ApIntOr_group_100",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 100
    -- shared split operator group (101) : OR_u32_u32_4027_inst 
    ApIntOr_group_101: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= iNsTr_252_4023 & iNsTr_249_4006;
      iNsTr_253_4028 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= OR_u32_u32_4027_inst_req_0;
      OR_u32_u32_4027_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= OR_u32_u32_4027_inst_req_1;
      OR_u32_u32_4027_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntOr",
          name => "ApIntOr_group_101",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 101
    -- shared split operator group (102) : SGT_f32_u1_2173_inst 
    ApFloatUgt_group_102: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= iNsTr_17_2155;
      iNsTr_25_2174 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= SGT_f32_u1_2173_inst_req_0;
      SGT_f32_u1_2173_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= SGT_f32_u1_2173_inst_req_1;
      SGT_f32_u1_2173_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApFloatUgt",
          name => "ApFloatUgt_group_102",
          input1_is_int => false, 
          input1_characteristic_width => 8, 
          input1_mantissa_width    => 23, 
          iwidth_1  => 32,
          input2_is_int => false, 
          input2_characteristic_width => 8, 
          input2_mantissa_width => 23, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "01000001111100000000000000000000",
          constant_width => 32,
          buffering  => 1,
          flow_through => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 102
    -- shared split operator group (103) : SGT_f32_u1_3615_inst 
    ApFloatUgt_group_103: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= iNsTr_85_3597;
      iNsTr_117_3616 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= SGT_f32_u1_3615_inst_req_0;
      SGT_f32_u1_3615_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= SGT_f32_u1_3615_inst_req_1;
      SGT_f32_u1_3615_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApFloatUgt",
          name => "ApFloatUgt_group_103",
          input1_is_int => false, 
          input1_characteristic_width => 8, 
          input1_mantissa_width    => 23, 
          iwidth_1  => 32,
          input2_is_int => false, 
          input2_characteristic_width => 8, 
          input2_mantissa_width => 23, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "01000010110010000000000000000000",
          constant_width => 32,
          buffering  => 1,
          flow_through => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 103
    -- shared split operator group (104) : SGT_f32_u1_3665_inst 
    ApFloatUgt_group_104: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= iNsTr_114_3647;
      iNsTr_151_3666 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= SGT_f32_u1_3665_inst_req_0;
      SGT_f32_u1_3665_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= SGT_f32_u1_3665_inst_req_1;
      SGT_f32_u1_3665_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApFloatUgt",
          name => "ApFloatUgt_group_104",
          input1_is_int => false, 
          input1_characteristic_width => 8, 
          input1_mantissa_width    => 23, 
          iwidth_1  => 32,
          input2_is_int => false, 
          input2_characteristic_width => 8, 
          input2_mantissa_width => 23, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "01000011010010000000000000000000",
          constant_width => 32,
          buffering  => 1,
          flow_through => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 104
    -- shared split operator group (105) : SGT_f64_u1_2123_inst 
    ApFloatUgt_group_105: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= iNsTr_13_2105;
      iNsTr_20_2124 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= SGT_f64_u1_2123_inst_req_0;
      SGT_f64_u1_2123_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= SGT_f64_u1_2123_inst_req_1;
      SGT_f64_u1_2123_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApFloatUgt",
          name => "ApFloatUgt_group_105",
          input1_is_int => false, 
          input1_characteristic_width => 11, 
          input1_mantissa_width    => 52, 
          iwidth_1  => 64,
          input2_is_int => false, 
          input2_characteristic_width => 11, 
          input2_mantissa_width => 52, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "0100000000101110000000000000000000000000000000000000000000000000",
          constant_width => 64,
          buffering  => 1,
          flow_through => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 105
    -- shared split operator group (106) : SGT_f64_u1_2209_inst 
    ApFloatUgt_group_106: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= iNsTr_22_2204;
      iNsTr_23_2210 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= SGT_f64_u1_2209_inst_req_0;
      SGT_f64_u1_2209_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= SGT_f64_u1_2209_inst_req_1;
      SGT_f64_u1_2209_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApFloatUgt",
          name => "ApFloatUgt_group_106",
          input1_is_int => false, 
          input1_characteristic_width => 11, 
          input1_mantissa_width    => 52, 
          iwidth_1  => 64,
          input2_is_int => false, 
          input2_characteristic_width => 11, 
          input2_mantissa_width => 52, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "0100000010011111010000000000000000000000000000000000000000000000",
          constant_width => 64,
          buffering  => 1,
          flow_through => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 106
    -- shared split operator group (107) : SGT_f64_u1_2222_inst 
    ApFloatUgt_group_107: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= iNsTr_22_2204;
      iNsTr_28_2223 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= SGT_f64_u1_2222_inst_req_0;
      SGT_f64_u1_2222_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= SGT_f64_u1_2222_inst_req_1;
      SGT_f64_u1_2222_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApFloatUgt",
          name => "ApFloatUgt_group_107",
          input1_is_int => false, 
          input1_characteristic_width => 11, 
          input1_mantissa_width    => 52, 
          iwidth_1  => 64,
          input2_is_int => false, 
          input2_characteristic_width => 11, 
          input2_mantissa_width => 52, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "0100000010100011100010000000000000000000000000000000000000000000",
          constant_width => 64,
          buffering  => 1,
          flow_through => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 107
    -- shared split operator group (108) : SGT_f64_u1_2255_inst 
    ApFloatUgt_group_108: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= iNsTr_22_2204;
      iNsTr_36_2256 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= SGT_f64_u1_2255_inst_req_0;
      SGT_f64_u1_2255_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= SGT_f64_u1_2255_inst_req_1;
      SGT_f64_u1_2255_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApFloatUgt",
          name => "ApFloatUgt_group_108",
          input1_is_int => false, 
          input1_characteristic_width => 11, 
          input1_mantissa_width    => 52, 
          iwidth_1  => 64,
          input2_is_int => false, 
          input2_characteristic_width => 11, 
          input2_mantissa_width => 52, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "0100000010100111011100000000000000000000000000000000000000000000",
          constant_width => 64,
          buffering  => 1,
          flow_through => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 108
    -- shared split operator group (109) : SHL_u32_u32_2354_inst 
    ApIntSHL_group_109: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= tmp10x_xix_xi30_2336;
      iNsTr_47_2355 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= SHL_u32_u32_2354_inst_req_0;
      SHL_u32_u32_2354_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= SHL_u32_u32_2354_inst_req_1;
      SHL_u32_u32_2354_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntSHL",
          name => "ApIntSHL_group_109",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000111",
          constant_width => 32,
          buffering  => 1,
          flow_through => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 109
    -- shared split operator group (110) : SHL_u32_u32_2424_inst 
    ApIntSHL_group_110: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= shifted_divisorx_x03x_xix_xix_xi34_2405;
      iNsTr_135_2425 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= SHL_u32_u32_2424_inst_req_0;
      SHL_u32_u32_2424_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= SHL_u32_u32_2424_inst_req_1;
      SHL_u32_u32_2424_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntSHL",
          name => "ApIntSHL_group_110",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000001",
          constant_width => 32,
          buffering  => 1,
          flow_through => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 110
    -- shared split operator group (111) : SHL_u32_u32_2430_inst 
    ApIntSHL_group_111: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= curr_quotientx_x02x_xix_xix_xi35_2412;
      iNsTr_136_2431 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= SHL_u32_u32_2430_inst_req_0;
      SHL_u32_u32_2430_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= SHL_u32_u32_2430_inst_req_1;
      SHL_u32_u32_2430_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntSHL",
          name => "ApIntSHL_group_111",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000001",
          constant_width => 32,
          buffering  => 1,
          flow_through => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 111
    -- shared split operator group (112) : SHL_u32_u32_2574_inst 
    ApIntSHL_group_112: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= tempx_x012x_xix_xi42_2563;
      iNsTr_206_2575 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= SHL_u32_u32_2574_inst_req_0;
      SHL_u32_u32_2574_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= SHL_u32_u32_2574_inst_req_1;
      SHL_u32_u32_2574_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntSHL",
          name => "ApIntSHL_group_112",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000001",
          constant_width => 32,
          buffering  => 1,
          flow_through => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 112
    -- shared split operator group (113) : SHL_u32_u32_2659_inst 
    ApIntSHL_group_113: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= expx_x0x_xlcssax_xix_xi49_2636;
      iNsTr_178_2660 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= SHL_u32_u32_2659_inst_req_0;
      SHL_u32_u32_2659_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= SHL_u32_u32_2659_inst_req_1;
      SHL_u32_u32_2659_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntSHL",
          name => "ApIntSHL_group_113",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000010111",
          constant_width => 32,
          buffering  => 1,
          flow_through => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 113
    -- shared split operator group (114) : SHL_u32_u32_2752_inst 
    ApIntSHL_group_114: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= tmp10x_xix_xi1_2706;
      iNsTr_68_2753 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= SHL_u32_u32_2752_inst_req_0;
      SHL_u32_u32_2752_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= SHL_u32_u32_2752_inst_req_1;
      SHL_u32_u32_2752_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntSHL",
          name => "ApIntSHL_group_114",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000111",
          constant_width => 32,
          buffering  => 1,
          flow_through => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 114
    -- shared split operator group (115) : SHL_u32_u32_2865_inst 
    ApIntSHL_group_115: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= shifted_divisorx_x03x_xix_xix_xi6_2847;
      iNsTr_199_2866 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= SHL_u32_u32_2865_inst_req_0;
      SHL_u32_u32_2865_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= SHL_u32_u32_2865_inst_req_1;
      SHL_u32_u32_2865_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntSHL",
          name => "ApIntSHL_group_115",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000001",
          constant_width => 32,
          buffering  => 1,
          flow_through => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 115
    -- shared split operator group (116) : SHL_u32_u32_2871_inst 
    ApIntSHL_group_116: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= curr_quotientx_x02x_xix_xix_xi7_2853;
      iNsTr_200_2872 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= SHL_u32_u32_2871_inst_req_0;
      SHL_u32_u32_2871_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= SHL_u32_u32_2871_inst_req_1;
      SHL_u32_u32_2871_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntSHL",
          name => "ApIntSHL_group_116",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000001",
          constant_width => 32,
          buffering  => 1,
          flow_through => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 116
    -- shared split operator group (117) : SHL_u32_u32_3008_inst 
    ApIntSHL_group_117: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= tempx_x012x_xix_xi17_2997;
      iNsTr_170_3009 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= SHL_u32_u32_3008_inst_req_0;
      SHL_u32_u32_3008_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= SHL_u32_u32_3008_inst_req_1;
      SHL_u32_u32_3008_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntSHL",
          name => "ApIntSHL_group_117",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000001",
          constant_width => 32,
          buffering  => 1,
          flow_through => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 117
    -- shared split operator group (118) : SHL_u32_u32_3098_inst 
    ApIntSHL_group_118: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= expx_x0x_xlcssax_xix_xi25_3075;
      iNsTr_130_3099 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= SHL_u32_u32_3098_inst_req_0;
      SHL_u32_u32_3098_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= SHL_u32_u32_3098_inst_req_1;
      SHL_u32_u32_3098_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntSHL",
          name => "ApIntSHL_group_118",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000010111",
          constant_width => 32,
          buffering  => 1,
          flow_through => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 118
    -- shared split operator group (119) : SHL_u32_u32_3198_inst 
    ApIntSHL_group_119: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= tmp10x_xix_xi_3145;
      iNsTr_92_3199 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= SHL_u32_u32_3198_inst_req_0;
      SHL_u32_u32_3198_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= SHL_u32_u32_3198_inst_req_1;
      SHL_u32_u32_3198_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntSHL",
          name => "ApIntSHL_group_119",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000111",
          constant_width => 32,
          buffering  => 1,
          flow_through => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 119
    -- shared split operator group (120) : SHL_u32_u32_3311_inst 
    ApIntSHL_group_120: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= shifted_divisorx_x03x_xix_xix_xi_3293;
      iNsTr_226_3312 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= SHL_u32_u32_3311_inst_req_0;
      SHL_u32_u32_3311_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= SHL_u32_u32_3311_inst_req_1;
      SHL_u32_u32_3311_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntSHL",
          name => "ApIntSHL_group_120",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000001",
          constant_width => 32,
          buffering  => 1,
          flow_through => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 120
    -- shared split operator group (121) : SHL_u32_u32_3317_inst 
    ApIntSHL_group_121: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= curr_quotientx_x02x_xix_xix_xi_3299;
      iNsTr_227_3318 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= SHL_u32_u32_3317_inst_req_0;
      SHL_u32_u32_3317_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= SHL_u32_u32_3317_inst_req_1;
      SHL_u32_u32_3317_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntSHL",
          name => "ApIntSHL_group_121",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000001",
          constant_width => 32,
          buffering  => 1,
          flow_through => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 121
    -- shared split operator group (122) : SHL_u32_u32_3454_inst 
    ApIntSHL_group_122: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= tempx_x012x_xix_xi_3443;
      iNsTr_194_3455 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= SHL_u32_u32_3454_inst_req_0;
      SHL_u32_u32_3454_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= SHL_u32_u32_3454_inst_req_1;
      SHL_u32_u32_3454_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntSHL",
          name => "ApIntSHL_group_122",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000001",
          constant_width => 32,
          buffering  => 1,
          flow_through => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 122
    -- shared split operator group (123) : SHL_u32_u32_3544_inst 
    ApIntSHL_group_123: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= expx_x0x_xlcssax_xix_xi_3521;
      iNsTr_159_3545 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= SHL_u32_u32_3544_inst_req_0;
      SHL_u32_u32_3544_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= SHL_u32_u32_3544_inst_req_1;
      SHL_u32_u32_3544_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntSHL",
          name => "ApIntSHL_group_123",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000010111",
          constant_width => 32,
          buffering  => 1,
          flow_through => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 123
    -- shared split operator group (124) : SHL_u32_u32_3706_inst 
    ApIntSHL_group_124: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= tmp10x_xi55_3701;
      iNsTr_147_3707 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= SHL_u32_u32_3706_inst_req_0;
      SHL_u32_u32_3706_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= SHL_u32_u32_3706_inst_req_1;
      SHL_u32_u32_3706_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntSHL",
          name => "ApIntSHL_group_124",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000111",
          constant_width => 32,
          buffering  => 1,
          flow_through => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 124
    -- shared split operator group (125) : SHL_u32_u32_3776_inst 
    ApIntSHL_group_125: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= shifted_divisorx_x03x_xix_xi_3757;
      iNsTr_234_3777 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= SHL_u32_u32_3776_inst_req_0;
      SHL_u32_u32_3776_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= SHL_u32_u32_3776_inst_req_1;
      SHL_u32_u32_3776_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntSHL",
          name => "ApIntSHL_group_125",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000001",
          constant_width => 32,
          buffering  => 1,
          flow_through => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 125
    -- shared split operator group (126) : SHL_u32_u32_3782_inst 
    ApIntSHL_group_126: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= curr_quotientx_x02x_xix_xi_3764;
      iNsTr_235_3783 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= SHL_u32_u32_3782_inst_req_0;
      SHL_u32_u32_3782_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= SHL_u32_u32_3782_inst_req_1;
      SHL_u32_u32_3782_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntSHL",
          name => "ApIntSHL_group_126",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000001",
          constant_width => 32,
          buffering  => 1,
          flow_through => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 126
    -- shared split operator group (127) : SHL_u32_u32_3926_inst 
    ApIntSHL_group_127: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= tempx_x012x_xi_3915;
      iNsTr_256_3927 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= SHL_u32_u32_3926_inst_req_0;
      SHL_u32_u32_3926_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= SHL_u32_u32_3926_inst_req_1;
      SHL_u32_u32_3926_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntSHL",
          name => "ApIntSHL_group_127",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000001",
          constant_width => 32,
          buffering  => 1,
          flow_through => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 127
    -- shared split operator group (128) : SHL_u32_u32_4011_inst 
    ApIntSHL_group_128: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= expx_x0x_xlcssax_xi_3988;
      iNsTr_250_4012 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= SHL_u32_u32_4011_inst_req_0;
      SHL_u32_u32_4011_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= SHL_u32_u32_4011_inst_req_1;
      SHL_u32_u32_4011_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntSHL",
          name => "ApIntSHL_group_128",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000010111",
          constant_width => 32,
          buffering  => 1,
          flow_through => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 128
    -- shared split operator group (129) : SLT_f32_u1_2160_inst 
    ApFloatUlt_group_129: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= iNsTr_17_2155;
      iNsTr_18_2161 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= SLT_f32_u1_2160_inst_req_0;
      SLT_f32_u1_2160_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= SLT_f32_u1_2160_inst_req_1;
      SLT_f32_u1_2160_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApFloatUlt",
          name => "ApFloatUlt_group_129",
          input1_is_int => false, 
          input1_characteristic_width => 8, 
          input1_mantissa_width    => 23, 
          iwidth_1  => 32,
          input2_is_int => false, 
          input2_characteristic_width => 8, 
          input2_mantissa_width => 23, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "11000001111100000000000000000000",
          constant_width => 32,
          buffering  => 1,
          flow_through => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 129
    -- shared split operator group (130) : SLT_f32_u1_3134_inst 
    ApFloatUlt_group_130: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= iNsTr_42_2683;
      iNsTr_60_3135 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= SLT_f32_u1_3134_inst_req_0;
      SLT_f32_u1_3134_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= SLT_f32_u1_3134_inst_req_1;
      SLT_f32_u1_3134_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApFloatUlt",
          name => "ApFloatUlt_group_130",
          input1_is_int => false, 
          input1_characteristic_width => 8, 
          input1_mantissa_width    => 23, 
          iwidth_1  => 32,
          input2_is_int => false, 
          input2_characteristic_width => 8, 
          input2_mantissa_width => 23, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "00111111100000000000000000000000",
          constant_width => 32,
          buffering  => 1,
          flow_through => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 130
    -- shared split operator group (131) : SLT_f32_u1_3602_inst 
    ApFloatUlt_group_131: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= iNsTr_85_3597;
      iNsTr_86_3603 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= SLT_f32_u1_3602_inst_req_0;
      SLT_f32_u1_3602_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= SLT_f32_u1_3602_inst_req_1;
      SLT_f32_u1_3602_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApFloatUlt",
          name => "ApFloatUlt_group_131",
          input1_is_int => false, 
          input1_characteristic_width => 8, 
          input1_mantissa_width    => 23, 
          iwidth_1  => 32,
          input2_is_int => false, 
          input2_characteristic_width => 8, 
          input2_mantissa_width => 23, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "11000010110010000000000000000000",
          constant_width => 32,
          buffering  => 1,
          flow_through => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 131
    -- shared split operator group (132) : SLT_f32_u1_3652_inst 
    ApFloatUlt_group_132: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= iNsTr_114_3647;
      iNsTr_115_3653 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= SLT_f32_u1_3652_inst_req_0;
      SLT_f32_u1_3652_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= SLT_f32_u1_3652_inst_req_1;
      SLT_f32_u1_3652_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApFloatUlt",
          name => "ApFloatUlt_group_132",
          input1_is_int => false, 
          input1_characteristic_width => 8, 
          input1_mantissa_width    => 23, 
          iwidth_1  => 32,
          input2_is_int => false, 
          input2_characteristic_width => 8, 
          input2_mantissa_width => 23, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "11000011010010000000000000000000",
          constant_width => 32,
          buffering  => 1,
          flow_through => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 132
    -- shared split operator group (133) : SLT_f64_u1_2110_inst 
    ApFloatUlt_group_133: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= iNsTr_13_2105;
      iNsTr_14_2111 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= SLT_f64_u1_2110_inst_req_0;
      SLT_f64_u1_2110_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= SLT_f64_u1_2110_inst_req_1;
      SLT_f64_u1_2110_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApFloatUlt",
          name => "ApFloatUlt_group_133",
          input1_is_int => false, 
          input1_characteristic_width => 11, 
          input1_mantissa_width    => 52, 
          iwidth_1  => 64,
          input2_is_int => false, 
          input2_characteristic_width => 11, 
          input2_mantissa_width => 52, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "1100000000101110000000000000000000000000000000000000000000000000",
          constant_width => 64,
          buffering  => 1,
          flow_through => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 133
    -- shared split operator group (134) : SUB_f32_f32_2082_inst SUB_f32_f32_3579_inst 
    ApFloatSub_group_134: Block -- 
      signal data_in: std_logic_vector(127 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 1, 1 => 1);
      -- 
    begin -- 
      data_in <= iNsTr_8_2078 & iNsTr_6_2075 & flux_refx_x0_2304 & iNsTr_42_2683;
      iNsTr_9_2083 <= data_out(63 downto 32);
      iNsTr_82_3580 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      reqL_unguarded(1) <= SUB_f32_f32_2082_inst_req_0;
      reqL_unguarded(0) <= SUB_f32_f32_3579_inst_req_0;
      SUB_f32_f32_2082_inst_ack_0 <= ackL_unguarded(1);
      SUB_f32_f32_3579_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= SUB_f32_f32_2082_inst_req_1;
      reqR_unguarded(0) <= SUB_f32_f32_3579_inst_req_1;
      SUB_f32_f32_2082_inst_ack_1 <= ackR_unguarded(1);
      SUB_f32_f32_3579_inst_ack_1 <= ackR_unguarded(0);
      ApFloatSub_group_134_accessRegulator_0: access_regulator_base generic map (name => "ApFloatSub_group_134_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      ApFloatSub_group_134_accessRegulator_1: access_regulator_base generic map (name => "ApFloatSub_group_134_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      gI: SplitGuardInterface generic map(nreqs => 2, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      PipedFpOp: PipelinedFPOperator -- 
        generic map( -- 
          name => "ApFloatSub_group_134",
          operator_id => "ApFloatSub",
          exponent_width => 8,
          fraction_width => 23, 
          no_arbitration => false,
          num_reqs => 2,
          use_input_buffering => true,
          detailed_buffering_per_input => inBUFs,
          detailed_buffering_per_output => outBUFs -- 
        )
        port map ( reqL => reqL , ackL => ackL, reqR => reqR, ackR => ackR, dataL => data_in, dataR => data_out, clk => clk, reset => reset); -- 
      -- 
    end Block; -- split operator group 134
    -- shared split operator group (135) : SUB_u32_u32_2478_inst 
    ApIntSub_group_135: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= xx_x016x_xix_xix_xi31_2370 & shifted_divisorx_x0x_xlcssax_xix_xix_xi37_2455;
      iNsTr_110_2479 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= SUB_u32_u32_2478_inst_req_0;
      SUB_u32_u32_2478_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= SUB_u32_u32_2478_inst_req_1;
      SUB_u32_u32_2478_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntSub",
          name => "ApIntSub_group_135",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 135
    -- shared split operator group (136) : SUB_u32_u32_2632_inst 
    ApIntSub_group_136: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= tmp25x_xix_xi46_2628 & xx_xlcssa15_2618;
      tmp26x_xix_xi47_2633 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= SUB_u32_u32_2632_inst_req_0;
      SUB_u32_u32_2632_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= SUB_u32_u32_2632_inst_req_1;
      SUB_u32_u32_2632_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntSub",
          name => "ApIntSub_group_136",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 136
    -- shared split operator group (137) : SUB_u32_u32_2798_inst 
    ApIntSub_group_137: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= iNsTr_65_2735 & iNsTr_67_2747;
      iNsTr_76_2799 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= SUB_u32_u32_2798_inst_req_0;
      SUB_u32_u32_2798_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= SUB_u32_u32_2798_inst_req_1;
      SUB_u32_u32_2798_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntSub",
          name => "ApIntSub_group_137",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 137
    -- shared split operator group (138) : SUB_u32_u32_2918_inst 
    ApIntSub_group_138: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= xx_x016x_xix_xix_xi3_2813 & shifted_divisorx_x0x_xlcssax_xix_xix_xi9_2896;
      iNsTr_166_2919 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= SUB_u32_u32_2918_inst_req_0;
      SUB_u32_u32_2918_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= SUB_u32_u32_2918_inst_req_1;
      SUB_u32_u32_2918_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntSub",
          name => "ApIntSub_group_138",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 138
    -- shared split operator group (139) : SUB_u32_u32_3066_inst 
    ApIntSub_group_139: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= tmp21x_xix_xi21_3062 & iNsTr_67_2747;
      tmp25x_xix_xi22_3067 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= SUB_u32_u32_3066_inst_req_0;
      SUB_u32_u32_3066_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= SUB_u32_u32_3066_inst_req_1;
      SUB_u32_u32_3066_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntSub",
          name => "ApIntSub_group_139",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 139
    -- shared split operator group (140) : SUB_u32_u32_3071_inst 
    ApIntSub_group_140: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= tmp25x_xix_xi22_3067 & xx_xlcssa10_3052;
      tmp26x_xix_xi23_3072 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= SUB_u32_u32_3071_inst_req_0;
      SUB_u32_u32_3071_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= SUB_u32_u32_3071_inst_req_1;
      SUB_u32_u32_3071_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntSub",
          name => "ApIntSub_group_140",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 140
    -- shared split operator group (141) : SUB_u32_u32_3244_inst 
    ApIntSub_group_141: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= iNsTr_89_3181 & iNsTr_91_3193;
      iNsTr_100_3245 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= SUB_u32_u32_3244_inst_req_0;
      SUB_u32_u32_3244_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= SUB_u32_u32_3244_inst_req_1;
      SUB_u32_u32_3244_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntSub",
          name => "ApIntSub_group_141",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 141
    -- shared split operator group (142) : SUB_u32_u32_3364_inst 
    ApIntSub_group_142: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= xx_x016x_xix_xix_xi_3259 & shifted_divisorx_x0x_xlcssax_xix_xix_xi_3342;
      iNsTr_190_3365 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= SUB_u32_u32_3364_inst_req_0;
      SUB_u32_u32_3364_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= SUB_u32_u32_3364_inst_req_1;
      SUB_u32_u32_3364_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntSub",
          name => "ApIntSub_group_142",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 142
    -- shared split operator group (143) : SUB_u32_u32_3512_inst 
    ApIntSub_group_143: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= tmp21x_xix_xi_3508 & iNsTr_91_3193;
      tmp25x_xix_xi_3513 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= SUB_u32_u32_3512_inst_req_0;
      SUB_u32_u32_3512_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= SUB_u32_u32_3512_inst_req_1;
      SUB_u32_u32_3512_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntSub",
          name => "ApIntSub_group_143",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 143
    -- shared split operator group (144) : SUB_u32_u32_3517_inst 
    ApIntSub_group_144: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= tmp25x_xix_xi_3513 & xx_xlcssa5_3498;
      tmp26x_xix_xi_3518 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= SUB_u32_u32_3517_inst_req_0;
      SUB_u32_u32_3517_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= SUB_u32_u32_3517_inst_req_1;
      SUB_u32_u32_3517_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntSub",
          name => "ApIntSub_group_144",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 144
    -- shared split operator group (145) : SUB_u32_u32_3830_inst 
    ApIntSub_group_145: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= xx_x016x_xix_xi_3722 & shifted_divisorx_x0x_xlcssax_xix_xi_3807;
      iNsTr_213_3831 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= SUB_u32_u32_3830_inst_req_0;
      SUB_u32_u32_3830_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= SUB_u32_u32_3830_inst_req_1;
      SUB_u32_u32_3830_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntSub",
          name => "ApIntSub_group_145",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 145
    -- shared split operator group (146) : SUB_u32_u32_3984_inst 
    ApIntSub_group_146: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= tmp25x_xi_3980 & xx_xlcssa_3970;
      tmp26x_xi_3985 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= SUB_u32_u32_3984_inst_req_0;
      SUB_u32_u32_3984_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= SUB_u32_u32_3984_inst_req_1;
      SUB_u32_u32_3984_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntSub",
          name => "ApIntSub_group_146",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 146
    -- shared split operator group (147) : UGT_u32_u1_2394_inst 
    ApIntUgt_group_147: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= iNsTr_78_2389;
      iNsTr_79_2395 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= UGT_u32_u1_2394_inst_req_0;
      UGT_u32_u1_2394_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= UGT_u32_u1_2394_inst_req_1;
      UGT_u32_u1_2394_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntUgt",
          name => "ApIntUgt_group_147",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "00000000000000011001111111100001",
          constant_width => 32,
          buffering  => 1,
          flow_through => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 147
    -- shared split operator group (148) : UGT_u32_u1_2836_inst 
    ApIntUgt_group_148: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= iNsTr_125_2832 & iNsTr_73_2783;
      iNsTr_126_2837 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= UGT_u32_u1_2836_inst_req_0;
      UGT_u32_u1_2836_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= UGT_u32_u1_2836_inst_req_1;
      UGT_u32_u1_2836_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntUgt",
          name => "ApIntUgt_group_148",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 148
    -- shared split operator group (149) : UGT_u32_u1_3282_inst 
    ApIntUgt_group_149: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= iNsTr_154_3278 & iNsTr_97_3229;
      iNsTr_155_3283 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= UGT_u32_u1_3282_inst_req_0;
      UGT_u32_u1_3282_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= UGT_u32_u1_3282_inst_req_1;
      UGT_u32_u1_3282_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntUgt",
          name => "ApIntUgt_group_149",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 149
    -- shared split operator group (150) : UGT_u32_u1_3746_inst 
    ApIntUgt_group_150: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= iNsTr_183_3741;
      iNsTr_184_3747 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= UGT_u32_u1_3746_inst_req_0;
      UGT_u32_u1_3746_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= UGT_u32_u1_3746_inst_req_1;
      UGT_u32_u1_3746_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntUgt",
          name => "ApIntUgt_group_150",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "00000000000000010100001111010111",
          constant_width => 32,
          buffering  => 1,
          flow_through => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 150
    -- shared split operator group (151) : ULT_u32_u1_2435_inst 
    ApIntUlt_group_151: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= iNsTr_135_2425 & iNsTr_78_2389;
      iNsTr_137_2436 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ULT_u32_u1_2435_inst_req_0;
      ULT_u32_u1_2435_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ULT_u32_u1_2435_inst_req_1;
      ULT_u32_u1_2435_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntUlt",
          name => "ApIntUlt_group_151",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 151
    -- shared split operator group (152) : ULT_u32_u1_2484_inst 
    ApIntUlt_group_152: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= iNsTr_110_2479;
      iNsTr_111_2485 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ULT_u32_u1_2484_inst_req_0;
      ULT_u32_u1_2484_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ULT_u32_u1_2484_inst_req_1;
      ULT_u32_u1_2484_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntUlt",
          name => "ApIntUlt_group_152",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "00000000000000011001111111100001",
          constant_width => 32,
          buffering  => 1,
          flow_through => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 152
    -- shared split operator group (153) : ULT_u32_u1_2876_inst 
    ApIntUlt_group_153: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= iNsTr_199_2866 & iNsTr_125_2832;
      iNsTr_201_2877 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ULT_u32_u1_2876_inst_req_0;
      ULT_u32_u1_2876_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ULT_u32_u1_2876_inst_req_1;
      ULT_u32_u1_2876_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntUlt",
          name => "ApIntUlt_group_153",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 153
    -- shared split operator group (154) : ULT_u32_u1_2923_inst 
    ApIntUlt_group_154: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= iNsTr_166_2919 & iNsTr_73_2783;
      iNsTr_167_2924 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ULT_u32_u1_2923_inst_req_0;
      ULT_u32_u1_2923_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ULT_u32_u1_2923_inst_req_1;
      ULT_u32_u1_2923_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntUlt",
          name => "ApIntUlt_group_154",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 154
    -- shared split operator group (155) : ULT_u32_u1_3322_inst 
    ApIntUlt_group_155: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= iNsTr_226_3312 & iNsTr_154_3278;
      iNsTr_228_3323 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ULT_u32_u1_3322_inst_req_0;
      ULT_u32_u1_3322_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ULT_u32_u1_3322_inst_req_1;
      ULT_u32_u1_3322_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntUlt",
          name => "ApIntUlt_group_155",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 155
    -- shared split operator group (156) : ULT_u32_u1_3369_inst 
    ApIntUlt_group_156: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= iNsTr_190_3365 & iNsTr_97_3229;
      iNsTr_191_3370 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ULT_u32_u1_3369_inst_req_0;
      ULT_u32_u1_3369_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ULT_u32_u1_3369_inst_req_1;
      ULT_u32_u1_3369_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntUlt",
          name => "ApIntUlt_group_156",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 156
    -- shared split operator group (157) : ULT_u32_u1_3787_inst 
    ApIntUlt_group_157: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= iNsTr_234_3777 & iNsTr_183_3741;
      iNsTr_236_3788 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ULT_u32_u1_3787_inst_req_0;
      ULT_u32_u1_3787_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ULT_u32_u1_3787_inst_req_1;
      ULT_u32_u1_3787_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntUlt",
          name => "ApIntUlt_group_157",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 157
    -- shared split operator group (158) : ULT_u32_u1_3836_inst 
    ApIntUlt_group_158: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= iNsTr_213_3831;
      iNsTr_214_3837 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ULT_u32_u1_3836_inst_req_0;
      ULT_u32_u1_3836_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ULT_u32_u1_3836_inst_req_1;
      ULT_u32_u1_3836_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntUlt",
          name => "ApIntUlt_group_158",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "00000000000000010100001111010111",
          constant_width => 32,
          buffering  => 1,
          flow_through => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 158
    -- shared split operator group (159) : XOR_u32_u32_2787_inst 
    ApIntXor_group_159: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= tmp6x_xix_xi2_2710 & tmp10x_xix_xi1_2706;
      iNsTr_74_2788 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= XOR_u32_u32_2787_inst_req_0;
      XOR_u32_u32_2787_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= XOR_u32_u32_2787_inst_req_1;
      XOR_u32_u32_2787_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntXor",
          name => "ApIntXor_group_159",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 159
    -- shared split operator group (160) : XOR_u32_u32_3233_inst 
    ApIntXor_group_160: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= tmp6x_xix_xi_3156 & tmp10x_xix_xi_3145;
      iNsTr_98_3234 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= XOR_u32_u32_3233_inst_req_0;
      XOR_u32_u32_3233_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= XOR_u32_u32_3233_inst_req_1;
      XOR_u32_u32_3233_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntXor",
          name => "ApIntXor_group_160",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 160
    -- shared split operator group (161) : switch_stmt_2800_select_expr_0 
    ApIntEq_group_161: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= iNsTr_73_2783;
      expr_2802_wire_constant_cmp <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= switch_stmt_2800_select_expr_0_req_0;
      switch_stmt_2800_select_expr_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= switch_stmt_2800_select_expr_0_req_1;
      switch_stmt_2800_select_expr_0_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntEq",
          name => "ApIntEq_group_161",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "00000000000000000000000000000000",
          constant_width => 32,
          buffering  => 1,
          flow_through => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 161
    -- shared split operator group (162) : switch_stmt_2800_select_expr_1 
    ApIntEq_group_162: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= iNsTr_73_2783;
      expr_2805_wire_constant_cmp <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= switch_stmt_2800_select_expr_1_req_0;
      switch_stmt_2800_select_expr_1_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= switch_stmt_2800_select_expr_1_req_1;
      switch_stmt_2800_select_expr_1_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntEq",
          name => "ApIntEq_group_162",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "00000000000000000000000000000001",
          constant_width => 32,
          buffering  => 1,
          flow_through => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 162
    -- shared split operator group (163) : switch_stmt_3246_select_expr_0 
    ApIntEq_group_163: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= iNsTr_97_3229;
      expr_3248_wire_constant_cmp <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= switch_stmt_3246_select_expr_0_req_0;
      switch_stmt_3246_select_expr_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= switch_stmt_3246_select_expr_0_req_1;
      switch_stmt_3246_select_expr_0_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntEq",
          name => "ApIntEq_group_163",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "00000000000000000000000000000000",
          constant_width => 32,
          buffering  => 1,
          flow_through => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 163
    -- shared split operator group (164) : switch_stmt_3246_select_expr_1 
    ApIntEq_group_164: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= iNsTr_97_3229;
      expr_3251_wire_constant_cmp <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= switch_stmt_3246_select_expr_1_req_0;
      switch_stmt_3246_select_expr_1_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= switch_stmt_3246_select_expr_1_req_1;
      switch_stmt_3246_select_expr_1_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntEq",
          name => "ApIntEq_group_164",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "00000000000000000000000000000001",
          constant_width => 32,
          buffering  => 1,
          flow_through => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 164
    -- shared split operator group (165) : type_cast_2104_inst 
    ApFloatResize_group_165: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= iNsTr_12_2100;
      iNsTr_13_2105 <= data_out(63 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= type_cast_2104_inst_req_0;
      type_cast_2104_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= type_cast_2104_inst_req_1;
      type_cast_2104_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApFloatResize",
          name => "ApFloatResize_group_165",
          input1_is_int => false, 
          input1_characteristic_width => 8, 
          input1_mantissa_width    => 23, 
          iwidth_1  => 32,
          input2_is_int => false, 
          input2_characteristic_width => 8, 
          input2_mantissa_width => 23, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => false,
          output_characteristic_width  => 11, 
          output_mantissa_width => 52, 
          owidth => 64,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 165
    -- shared split operator group (166) : type_cast_2203_inst 
    ApFloatResize_group_166: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= iNsTr_8_2078;
      iNsTr_22_2204 <= data_out(63 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= type_cast_2203_inst_req_0;
      type_cast_2203_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= type_cast_2203_inst_req_1;
      type_cast_2203_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApFloatResize",
          name => "ApFloatResize_group_166",
          input1_is_int => false, 
          input1_characteristic_width => 8, 
          input1_mantissa_width    => 23, 
          iwidth_1  => 32,
          input2_is_int => false, 
          input2_characteristic_width => 8, 
          input2_mantissa_width => 23, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => false,
          output_characteristic_width  => 11, 
          output_mantissa_width => 52, 
          owidth => 64,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 166
    -- shared split operator group (167) : type_cast_2536_inst 
    ApIntToApIntSigned_group_167: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= xx_xlcssa19_2493;
      type_cast_2536_wire <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= type_cast_2536_inst_req_0;
      type_cast_2536_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= type_cast_2536_inst_req_1;
      type_cast_2536_inst_ack_1 <= ackR_unguarded(0);
      reqL <= reqL_unguarded;
      reqR <= reqR_unguarded;
      ackL_unguarded <= ackL;
      ackR_unguarded <= ackR;
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntToApIntSigned",
          name => "ApIntToApIntSigned_group_167",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => true,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 167
    -- shared split operator group (168) : type_cast_2590_inst 
    ApIntToApIntSigned_group_168: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= iNsTr_206_2575;
      type_cast_2590_wire <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= type_cast_2590_inst_req_0;
      type_cast_2590_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= type_cast_2590_inst_req_1;
      type_cast_2590_inst_ack_1 <= ackR_unguarded(0);
      reqL <= reqL_unguarded;
      reqR <= reqR_unguarded;
      ackL_unguarded <= ackL;
      ackR_unguarded <= ackR;
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntToApIntSigned",
          name => "ApIntToApIntSigned_group_168",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => true,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 168
    -- shared split operator group (169) : type_cast_2970_inst 
    ApIntToApIntSigned_group_169: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= tempx_x0x_xphx_xix_xi14_2949;
      type_cast_2970_wire <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= type_cast_2970_inst_req_0;
      type_cast_2970_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= type_cast_2970_inst_req_1;
      type_cast_2970_inst_ack_1 <= ackR_unguarded(0);
      reqL <= reqL_unguarded;
      reqR <= reqR_unguarded;
      ackL_unguarded <= ackL;
      ackR_unguarded <= ackR;
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntToApIntSigned",
          name => "ApIntToApIntSigned_group_169",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => true,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 169
    -- shared split operator group (170) : type_cast_3024_inst 
    ApIntToApIntSigned_group_170: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= iNsTr_170_3009;
      type_cast_3024_wire <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= type_cast_3024_inst_req_0;
      type_cast_3024_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= type_cast_3024_inst_req_1;
      type_cast_3024_inst_ack_1 <= ackR_unguarded(0);
      reqL <= reqL_unguarded;
      reqR <= reqR_unguarded;
      ackL_unguarded <= ackL;
      ackR_unguarded <= ackR;
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntToApIntSigned",
          name => "ApIntToApIntSigned_group_170",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => true,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 170
    -- shared split operator group (171) : type_cast_3416_inst 
    ApIntToApIntSigned_group_171: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= tempx_x0x_xphx_xix_xi_3395;
      type_cast_3416_wire <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= type_cast_3416_inst_req_0;
      type_cast_3416_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= type_cast_3416_inst_req_1;
      type_cast_3416_inst_ack_1 <= ackR_unguarded(0);
      reqL <= reqL_unguarded;
      reqR <= reqR_unguarded;
      ackL_unguarded <= ackL;
      ackR_unguarded <= ackR;
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntToApIntSigned",
          name => "ApIntToApIntSigned_group_171",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => true,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 171
    -- shared split operator group (172) : type_cast_3470_inst 
    ApIntToApIntSigned_group_172: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= iNsTr_194_3455;
      type_cast_3470_wire <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= type_cast_3470_inst_req_0;
      type_cast_3470_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= type_cast_3470_inst_req_1;
      type_cast_3470_inst_ack_1 <= ackR_unguarded(0);
      reqL <= reqL_unguarded;
      reqR <= reqR_unguarded;
      ackL_unguarded <= ackL;
      ackR_unguarded <= ackR;
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntToApIntSigned",
          name => "ApIntToApIntSigned_group_172",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => true,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 172
    -- shared split operator group (173) : type_cast_3888_inst 
    ApIntToApIntSigned_group_173: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= xx_xlcssa4_3845;
      type_cast_3888_wire <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= type_cast_3888_inst_req_0;
      type_cast_3888_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= type_cast_3888_inst_req_1;
      type_cast_3888_inst_ack_1 <= ackR_unguarded(0);
      reqL <= reqL_unguarded;
      reqR <= reqR_unguarded;
      ackL_unguarded <= ackL;
      ackR_unguarded <= ackR;
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntToApIntSigned",
          name => "ApIntToApIntSigned_group_173",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => true,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 173
    -- shared split operator group (174) : type_cast_3942_inst 
    ApIntToApIntSigned_group_174: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= iNsTr_256_3927;
      type_cast_3942_wire <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= type_cast_3942_inst_req_0;
      type_cast_3942_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= type_cast_3942_inst_req_1;
      type_cast_3942_inst_ack_1 <= ackR_unguarded(0);
      reqL <= reqL_unguarded;
      reqR <= reqR_unguarded;
      ackL_unguarded <= ackL;
      ackR_unguarded <= ackR;
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntToApIntSigned",
          name => "ApIntToApIntSigned_group_174",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => true,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 174
    -- shared inport operator group (0) : RPIPE_in_data_2071_inst RPIPE_in_data_2077_inst RPIPE_in_data_2068_inst RPIPE_in_data_2074_inst 
    InportGroup0: Block -- 
      signal data_out: std_logic_vector(127 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 3 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 3 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 3 downto 0);
      signal guard_vector : std_logic_vector( 3 downto 0);
      constant outBUFs : IntegerArray(3 downto 0) := (3 => 1, 2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(3 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false);
      constant guardBuffering: IntegerArray(3 downto 0)  := (0 => 1, 1 => 1, 2 => 1, 3 => 1);
      -- 
    begin -- 
      reqL_unguarded(3) <= RPIPE_in_data_2071_inst_req_0;
      reqL_unguarded(2) <= RPIPE_in_data_2077_inst_req_0;
      reqL_unguarded(1) <= RPIPE_in_data_2068_inst_req_0;
      reqL_unguarded(0) <= RPIPE_in_data_2074_inst_req_0;
      RPIPE_in_data_2071_inst_ack_0 <= ackL_unguarded(3);
      RPIPE_in_data_2077_inst_ack_0 <= ackL_unguarded(2);
      RPIPE_in_data_2068_inst_ack_0 <= ackL_unguarded(1);
      RPIPE_in_data_2074_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(3) <= RPIPE_in_data_2071_inst_req_1;
      reqR_unguarded(2) <= RPIPE_in_data_2077_inst_req_1;
      reqR_unguarded(1) <= RPIPE_in_data_2068_inst_req_1;
      reqR_unguarded(0) <= RPIPE_in_data_2074_inst_req_1;
      RPIPE_in_data_2071_inst_ack_1 <= ackR_unguarded(3);
      RPIPE_in_data_2077_inst_ack_1 <= ackR_unguarded(2);
      RPIPE_in_data_2068_inst_ack_1 <= ackR_unguarded(1);
      RPIPE_in_data_2074_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      gI: SplitGuardInterface generic map(nreqs => 4, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      iNsTr_4_2072 <= data_out(127 downto 96);
      iNsTr_8_2078 <= data_out(95 downto 64);
      iNsTr_2_2069 <= data_out(63 downto 32);
      iNsTr_6_2075 <= data_out(31 downto 0);
      in_data_read_0: InputPortFullRate -- 
        generic map ( name => "in_data_read_0", data_width => 32,  num_reqs => 4,  output_buffering => outBUFs,   no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => in_data_pipe_read_req(0),
          oack => in_data_pipe_read_ack(0),
          odata => in_data_pipe_read_data(31 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared outport operator group (0) : WPIPE_out_data_4043_inst WPIPE_out_data_4046_inst WPIPE_out_data_4049_inst WPIPE_out_data_4052_inst 
    OutportGroup0: Block -- 
      signal data_in: std_logic_vector(127 downto 0);
      signal sample_req, sample_ack : BooleanArray( 3 downto 0);
      signal update_req, update_ack : BooleanArray( 3 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 3 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 3 downto 0);
      signal guard_vector : std_logic_vector( 3 downto 0);
      constant inBUFs : IntegerArray(3 downto 0) := (3 => 1, 2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(3 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false);
      constant guardBuffering: IntegerArray(3 downto 0)  := (0 => 1, 1 => 1, 2 => 1, 3 => 1);
      -- 
    begin -- 
      sample_req_unguarded(3) <= WPIPE_out_data_4043_inst_req_0;
      sample_req_unguarded(2) <= WPIPE_out_data_4046_inst_req_0;
      sample_req_unguarded(1) <= WPIPE_out_data_4049_inst_req_0;
      sample_req_unguarded(0) <= WPIPE_out_data_4052_inst_req_0;
      WPIPE_out_data_4043_inst_ack_0 <= sample_ack_unguarded(3);
      WPIPE_out_data_4046_inst_ack_0 <= sample_ack_unguarded(2);
      WPIPE_out_data_4049_inst_ack_0 <= sample_ack_unguarded(1);
      WPIPE_out_data_4052_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(3) <= WPIPE_out_data_4043_inst_req_1;
      update_req_unguarded(2) <= WPIPE_out_data_4046_inst_req_1;
      update_req_unguarded(1) <= WPIPE_out_data_4049_inst_req_1;
      update_req_unguarded(0) <= WPIPE_out_data_4052_inst_req_1;
      WPIPE_out_data_4043_inst_ack_1 <= update_ack_unguarded(3);
      WPIPE_out_data_4046_inst_ack_1 <= update_ack_unguarded(2);
      WPIPE_out_data_4049_inst_ack_1 <= update_ack_unguarded(1);
      WPIPE_out_data_4052_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      gI: SplitGuardInterface generic map(nreqs => 4, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      data_in <= iNsTr_216_4035 & iNsTr_81_3568 & iNsTr_59_3122 & iNsTr_42_2683;
      out_data_write_0: OutputPortFullRate -- 
        generic map ( name => "out_data", data_width => 32, num_reqs => 4, input_buffering => inBUFs, no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => out_data_pipe_write_req(0),
          oack => out_data_pipe_write_ack(0),
          odata => out_data_pipe_write_data(31 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- 
  end Block; -- data_path
  -- 
end Default;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;
library work;
use work.ahir_system_global_package.all;
entity ahir_system is  -- system 
  port (-- 
    clk : in std_logic;
    reset : in std_logic;
    in_data_pipe_write_data: in std_logic_vector(31 downto 0);
    in_data_pipe_write_req : in std_logic_vector(0 downto 0);
    in_data_pipe_write_ack : out std_logic_vector(0 downto 0);
    out_data_pipe_read_data: out std_logic_vector(31 downto 0);
    out_data_pipe_read_req : in std_logic_vector(0 downto 0);
    out_data_pipe_read_ack : out std_logic_vector(0 downto 0)); -- 
  -- 
end entity; 
architecture Default of ahir_system is -- system-architecture 
  -- declarations related to module vector_control_daemon
  component vector_control_daemon is -- 
    generic (tag_length : integer); 
    port ( -- 
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic;
      in_data_pipe_read_req : out  std_logic_vector(0 downto 0);
      in_data_pipe_read_ack : in   std_logic_vector(0 downto 0);
      in_data_pipe_read_data : in   std_logic_vector(31 downto 0);
      out_data_pipe_write_req : out  std_logic_vector(0 downto 0);
      out_data_pipe_write_ack : in   std_logic_vector(0 downto 0);
      out_data_pipe_write_data : out  std_logic_vector(31 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) -- 
    );
    -- 
  end component;
  -- argument signals for module vector_control_daemon
  signal vector_control_daemon_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal vector_control_daemon_tag_out   : std_logic_vector(1 downto 0);
  signal vector_control_daemon_start_req : std_logic;
  signal vector_control_daemon_start_ack : std_logic;
  signal vector_control_daemon_fin_req   : std_logic;
  signal vector_control_daemon_fin_ack : std_logic;
  -- aggregate signals for read from pipe in_data
  signal in_data_pipe_read_data: std_logic_vector(31 downto 0);
  signal in_data_pipe_read_req: std_logic_vector(0 downto 0);
  signal in_data_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe out_data
  signal out_data_pipe_write_data: std_logic_vector(31 downto 0);
  signal out_data_pipe_write_req: std_logic_vector(0 downto 0);
  signal out_data_pipe_write_ack: std_logic_vector(0 downto 0);
  -- 
begin -- 
  -- module vector_control_daemon
  vector_control_daemon_instance:vector_control_daemon-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => vector_control_daemon_start_req,
      start_ack => vector_control_daemon_start_ack,
      fin_req => vector_control_daemon_fin_req,
      fin_ack => vector_control_daemon_fin_ack,
      clk => clk,
      reset => reset,
      in_data_pipe_read_req => in_data_pipe_read_req(0 downto 0),
      in_data_pipe_read_ack => in_data_pipe_read_ack(0 downto 0),
      in_data_pipe_read_data => in_data_pipe_read_data(31 downto 0),
      out_data_pipe_write_req => out_data_pipe_write_req(0 downto 0),
      out_data_pipe_write_ack => out_data_pipe_write_ack(0 downto 0),
      out_data_pipe_write_data => out_data_pipe_write_data(31 downto 0),
      tag_in => vector_control_daemon_tag_in,
      tag_out => vector_control_daemon_tag_out-- 
    ); -- 
  -- module will be run forever 
  vector_control_daemon_tag_in <= (others => '0');
  vector_control_daemon_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => vector_control_daemon_start_req, start_ack => vector_control_daemon_start_ack,  fin_req => vector_control_daemon_fin_req,  fin_ack => vector_control_daemon_fin_ack);
  in_data_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe in_data",
      num_reads => 1,
      num_writes => 1,
      data_width => 32,
      lifo_mode => false,
      depth => 1 --
    )
    port map( -- 
      read_req => in_data_pipe_read_req,
      read_ack => in_data_pipe_read_ack,
      read_data => in_data_pipe_read_data,
      write_req => in_data_pipe_write_req,
      write_ack => in_data_pipe_write_ack,
      write_data => in_data_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  out_data_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe out_data",
      num_reads => 1,
      num_writes => 1,
      data_width => 32,
      lifo_mode => false,
      depth => 1 --
    )
    port map( -- 
      read_req => out_data_pipe_read_req,
      read_ack => out_data_pipe_read_ack,
      read_data => out_data_pipe_read_data,
      write_req => out_data_pipe_write_req,
      write_ack => out_data_pipe_write_ack,
      write_data => out_data_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  -- 
end Default;
